* SPICE3 file created from carry_select_adder.ext - technology: sky130A

V17 cin0 GND 0
V18 cin1 GND 1.8
vdd vdd GND 1.8
V1 a0 GND PULSE(1.8 0 0 .1n .1n 80 90n 1)
V2 a1 GND PULSE(1.8 0 0 .1n .1n 40n 80n 2)
V3 a2 GND PULSE(1.8 0 0 .1n .1n 20n 40n 3)
V4 a3 GND PULSE(1.8 0 0 .1n .1n 10n 20n 4)
V5 a4 GND PULSE(0 1.8 0 .1n .1n 80 90n 1)
V6 a5 GND PULSE(0 1.8 0 .1n .1n 40n 80n 2)
V7 a6 GND PULSE(0 1.8 0 .1n .1n 20n 40n 3)
V8 a7 GND PULSE(0 1.8 0 .1n .1n 10n 20n 4)
V9 b0 GND PULSE(1.8 0 0 .1n .1n 80 90n 1)
V10 b1 GND PULSE(1.8 0 0 .1n .1n 40n 80n 2)
V11 b2 GND PULSE(1.8 0 0 .1n .1n 20n 40n 3)
V12 b3 GND PULSE(1.8 0 0 .1n .1n 10n 20n 4)
V13 b4 GND PULSE(0 1.8 0 .1n .1n 80 90n 1)
V14 b5 GND PULSE(0 1.8 0 .1n .1n 40n 80n 2)
V15 b6 GND PULSE(0 1.8 0 .1n .1n 20n 40n 3)
V16 b7 GND PULSE(0 1.8 0 .1n .1n 10n 20n 4)


.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.tran .02ns 80ns
.save all


X0 full_adder_10/a_760_n530# b6 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.315 pd=2.5 as=0.315 ps=2.5 w=0.9 l=0.15
X1 full_adder_10/a_510_n530# a6 full_adder_10/a_760_n530# gnd sky130_fd_pr__nfet_01v8 ad=0.315 pd=2.5 as=0.315 ps=2.5 w=0.9 l=0.15
X2 full_adder_11/cin full_adder_10/a_510_n530# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0.315 ps=2.5 w=0.9 l=0.15
X3 full_adder_10/a_10_40# b6 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.63 pd=4.3 as=0.63 ps=4.3 w=1.8 l=0.15
X4 full_adder_10/a_1260_40# full_adder_8/cout vdd vdd sky130_fd_pr__pfet_01v8 ad=0.63 pd=4.3 as=0.63 ps=4.3 w=1.8 l=0.15
X5 full_adder_10/a_2260_40# a6 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.63 pd=4.3 as=0.63 ps=4.3 w=1.8 l=0.15
X6 full_adder_10/a_10_n530# b6 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.315 pd=2.5 as=0.315 ps=2.5 w=0.9 l=0.15
X7 full_adder_10/a_510_n530# full_adder_8/cout full_adder_10/a_10_n530# gnd sky130_fd_pr__nfet_01v8 ad=0.315 pd=2.5 as=0.315 ps=2.5 w=0.9 l=0.15
X8 full_adder_11/cin full_adder_10/a_510_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0.1575 ps=1.6 w=0.45 l=0.15
X9 full_adder_10/a_510_n530# a6 full_adder_10/a_760_40# vdd sky130_fd_pr__pfet_01v8 ad=0.63 pd=4.3 as=0.63 ps=4.3 w=1.8 l=0.15
X10 mux_2to1_2/in2 full_adder_10/a_2010_n530# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0.315 ps=2.5 w=0.9 l=0.15
X11 full_adder_10/a_2010_n530# full_adder_10/a_2670_n140# full_adder_10/a_2510_n530# gnd sky130_fd_pr__nfet_01v8 ad=0.315 pd=2.5 as=0.315 ps=2.5 w=0.9 l=0.15
X12 mux_2to1_2/in2 full_adder_10/a_2010_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0.1575 ps=1.6 w=0.45 l=0.15
X13 full_adder_10/a_1260_40# a6 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.63 pd=4.3 as=0.63 ps=4.3 w=1.8 l=0.15
X14 full_adder_10/a_510_n530# full_adder_8/cout full_adder_10/a_10_40# vdd sky130_fd_pr__pfet_01v8 ad=0.63 pd=4.3 as=0.63 ps=4.3 w=1.8 l=0.15
X15 full_adder_10/a_1260_n530# full_adder_8/cout gnd gnd sky130_fd_pr__nfet_01v8 ad=0.315 pd=2.5 as=0.315 ps=2.5 w=0.9 l=0.15
X16 full_adder_10/a_2010_n530# full_adder_10/a_510_n530# full_adder_10/a_1260_n530# gnd sky130_fd_pr__nfet_01v8 ad=0.315 pd=2.5 as=0.315 ps=2.5 w=0.9 l=0.15
X17 full_adder_10/a_2510_40# b6 full_adder_10/a_2260_40# vdd sky130_fd_pr__pfet_01v8 ad=0.63 pd=4.3 as=0.63 ps=4.3 w=1.8 l=0.15
X18 full_adder_10/a_2010_n530# full_adder_10/a_510_n530# full_adder_10/a_1260_40# vdd sky130_fd_pr__pfet_01v8 ad=0.63 pd=4.3 as=0.63 ps=4.3 w=1.8 l=0.15
X19 full_adder_10/a_2260_n530# a6 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.315 pd=2.5 as=0.315 ps=2.5 w=0.9 l=0.15
X20 full_adder_10/a_2510_n530# b6 full_adder_10/a_2260_n530# gnd sky130_fd_pr__nfet_01v8 ad=0.315 pd=2.5 as=0.315 ps=2.5 w=0.9 l=0.15
X21 full_adder_10/a_10_n530# a6 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.315 pd=2.5 as=0.315 ps=2.5 w=0.9 l=0.15
X22 full_adder_10/a_10_40# a6 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.63 pd=4.3 as=0.63 ps=4.3 w=1.8 l=0.15
X23 full_adder_10/a_1260_n530# a6 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.315 pd=2.5 as=0.315 ps=2.5 w=0.9 l=0.15
X24 full_adder_10/a_1260_n530# b6 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.315 pd=2.5 as=0.315 ps=2.5 w=0.9 l=0.15
X25 full_adder_10/a_760_40# b6 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.63 pd=4.3 as=0.63 ps=4.3 w=1.8 l=0.15
X26 full_adder_10/a_1260_40# b6 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.63 pd=4.3 as=0.63 ps=4.3 w=1.8 l=0.15
X27 full_adder_10/a_2010_n530# full_adder_10/a_2670_n140# full_adder_10/a_2510_40# vdd sky130_fd_pr__pfet_01v8 ad=0.63 pd=4.3 as=0.63 ps=4.3 w=1.8 l=0.15
X28 full_adder_11/a_760_n530# b7 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=31.0275 ps=256.4 w=0.9 l=0.15
X29 full_adder_11/a_510_n530# a7 full_adder_11/a_760_n530# gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X30 mux_2to1_4/in2 full_adder_11/a_510_n530# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.4725 pd=4.1 as=56.7 ps=396.1 w=0.9 l=0.15
X31 full_adder_11/a_10_40# b7 vdd vdd sky130_fd_pr__pfet_01v8 ad=1.89 pd=12.9 as=0 ps=0 w=1.8 l=0.15
X32 full_adder_11/a_1260_40# full_adder_11/cin vdd vdd sky130_fd_pr__pfet_01v8 ad=2.52 pd=17.2 as=0 ps=0 w=1.8 l=0.15
X33 full_adder_11/a_2260_40# a7 vdd vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=0 ps=0 w=1.8 l=0.15
X34 full_adder_11/a_10_n530# b7 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.945 pd=7.5 as=0 ps=0 w=0.9 l=0.15
X35 full_adder_11/a_510_n530# full_adder_11/cin full_adder_11/a_10_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X36 mux_2to1_4/in2 full_adder_11/a_510_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.315 pd=3.2 as=0 ps=0 w=0.45 l=0.15
X37 full_adder_11/a_510_n530# a7 full_adder_11/a_760_40# vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=1.26 ps=8.6 w=1.8 l=0.15
X38 mux_2to1_3/in2 full_adder_11/a_2010_n530# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.4725 pd=4.1 as=0 ps=0 w=0.9 l=0.15
X39 full_adder_11/a_2010_n530# full_adder_11/a_2670_n140# full_adder_11/a_2510_n530# gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0.63 ps=5 w=0.9 l=0.15
X40 mux_2to1_3/in2 full_adder_11/a_2010_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.315 pd=3.2 as=0 ps=0 w=0.45 l=0.15
X41 full_adder_11/a_1260_40# a7 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X42 full_adder_11/a_510_n530# full_adder_11/cin full_adder_11/a_10_40# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X43 full_adder_11/a_1260_n530# full_adder_11/cin gnd gnd sky130_fd_pr__nfet_01v8 ad=1.26 pd=10 as=0 ps=0 w=0.9 l=0.15
X44 full_adder_11/a_2010_n530# full_adder_11/a_510_n530# full_adder_11/a_1260_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X45 full_adder_11/a_2510_40# b7 full_adder_11/a_2260_40# vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=0 ps=0 w=1.8 l=0.15
X46 full_adder_11/a_2010_n530# full_adder_11/a_510_n530# full_adder_11/a_1260_40# vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=0 ps=0 w=1.8 l=0.15
X47 full_adder_11/a_2260_n530# a7 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X48 full_adder_11/a_2510_n530# b7 full_adder_11/a_2260_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X49 full_adder_11/a_10_n530# a7 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X50 full_adder_11/a_10_40# a7 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X51 full_adder_11/a_1260_n530# a7 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X52 full_adder_11/a_1260_n530# b7 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X53 full_adder_11/a_760_40# b7 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X54 full_adder_11/a_1260_40# b7 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X55 full_adder_11/a_2010_n530# full_adder_11/a_2670_n140# full_adder_11/a_2510_40# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X56 s4 mux_2to1_0/a_2510_640# mux_2to1_0/in1 gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0.1575 ps=1.6 w=0.45 l=0.15
X57 s4 mux_2to1_4/sel mux_2to1_0/in2 gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0.1575 ps=1.6 w=0.45 l=0.15
X58 mux_2to1_0/a_2510_640# mux_2to1_4/sel gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0.1575 ps=1.6 w=0.45 l=0.15
X59 s4 mux_2to1_4/sel mux_2to1_0/in1 mux_2to1_0/vdd sky130_fd_pr__pfet_01v8 ad=0.1575 pd=1.6 as=0.1575 ps=1.6 w=0.45 l=0.15
X60 s4 mux_2to1_0/a_2510_640# mux_2to1_0/in2 mux_2to1_0/vdd sky130_fd_pr__pfet_01v8 ad=0.1575 pd=1.6 as=0.1575 ps=1.6 w=0.45 l=0.15
X61 mux_2to1_0/a_2510_640# mux_2to1_4/sel mux_2to1_0/vdd mux_2to1_0/vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0.315 ps=2.5 w=0.9 l=0.15
X62 s5 mux_2to1_1/a_2510_640# mux_2to1_1/in1 gnd sky130_fd_pr__nfet_01v8 ad=0.315 pd=3.2 as=0.315 ps=3.2 w=0.45 l=0.15
X63 s5 mux_2to1_4/sel mux_2to1_1/in2 gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.315 ps=3.2 w=0.45 l=0.15
X64 mux_2to1_1/a_2510_640# mux_2to1_4/sel gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X65 s5 mux_2to1_4/sel mux_2to1_1/in1 vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=3.2 as=0.4725 ps=4.1 w=0.45 l=0.15
X66 s5 mux_2to1_1/a_2510_640# mux_2to1_1/in2 vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.4725 ps=4.1 w=0.45 l=0.15
X67 mux_2to1_1/a_2510_640# mux_2to1_4/sel vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X68 s6 mux_2to1_2/a_2510_640# mux_2to1_2/in1 gnd sky130_fd_pr__nfet_01v8 ad=0.315 pd=3.2 as=0.315 ps=3.2 w=0.45 l=0.15
X69 s6 mux_2to1_4/sel mux_2to1_2/in2 gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.315 ps=3.2 w=0.45 l=0.15
X70 mux_2to1_2/a_2510_640# mux_2to1_4/sel gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X71 s6 mux_2to1_4/sel mux_2to1_2/in1 vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=3.2 as=0.4725 ps=4.1 w=0.45 l=0.15
X72 s6 mux_2to1_2/a_2510_640# mux_2to1_2/in2 vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.4725 ps=4.1 w=0.45 l=0.15
X73 mux_2to1_2/a_2510_640# mux_2to1_4/sel vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X74 s7 mux_2to1_3/a_2510_640# mux_2to1_3/in1 gnd sky130_fd_pr__nfet_01v8 ad=0.315 pd=3.2 as=0.315 ps=3.2 w=0.45 l=0.15
X75 s7 mux_2to1_4/sel mux_2to1_3/in2 gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.45 l=0.15
X76 mux_2to1_3/a_2510_640# mux_2to1_4/sel gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X77 s7 mux_2to1_4/sel mux_2to1_3/in1 vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=3.2 as=0.4725 ps=4.1 w=0.45 l=0.15
X78 s7 mux_2to1_3/a_2510_640# mux_2to1_3/in2 vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.45 l=0.15
X79 mux_2to1_3/a_2510_640# mux_2to1_4/sel vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X80 full_adder_0/a_760_n530# b1 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X81 full_adder_0/a_510_n530# a1 full_adder_0/a_760_n530# gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X82 full_adder_2/cin full_adder_0/a_510_n530# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X83 full_adder_0/a_10_40# b1 vdd vdd sky130_fd_pr__pfet_01v8 ad=1.89 pd=12.9 as=0 ps=0 w=1.8 l=0.15
X84 full_adder_0/a_1260_40# full_adder_0/cin vdd vdd sky130_fd_pr__pfet_01v8 ad=2.52 pd=17.2 as=0 ps=0 w=1.8 l=0.15
X85 full_adder_0/a_2260_40# a1 vdd vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=0 ps=0 w=1.8 l=0.15
X86 full_adder_0/a_10_n530# b1 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.945 pd=7.5 as=0 ps=0 w=0.9 l=0.15
X87 full_adder_0/a_510_n530# full_adder_0/cin full_adder_0/a_10_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X88 full_adder_2/cin full_adder_0/a_510_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X89 full_adder_0/a_510_n530# a1 full_adder_0/a_760_40# vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=1.26 ps=8.6 w=1.8 l=0.15
X90 s1 full_adder_0/a_2010_n530# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X91 full_adder_0/a_2010_n530# full_adder_0/a_2670_n140# full_adder_0/a_2510_n530# gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0.63 ps=5 w=0.9 l=0.15
X92 s1 full_adder_0/a_2010_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X93 full_adder_0/a_1260_40# a1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X94 full_adder_0/a_510_n530# full_adder_0/cin full_adder_0/a_10_40# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X95 full_adder_0/a_1260_n530# full_adder_0/cin gnd gnd sky130_fd_pr__nfet_01v8 ad=1.26 pd=10 as=0 ps=0 w=0.9 l=0.15
X96 full_adder_0/a_2010_n530# full_adder_0/a_510_n530# full_adder_0/a_1260_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X97 full_adder_0/a_2510_40# b1 full_adder_0/a_2260_40# vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=0 ps=0 w=1.8 l=0.15
X98 full_adder_0/a_2010_n530# full_adder_0/a_510_n530# full_adder_0/a_1260_40# vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=0 ps=0 w=1.8 l=0.15
X99 full_adder_0/a_2260_n530# a1 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X100 full_adder_0/a_2510_n530# b1 full_adder_0/a_2260_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X101 full_adder_0/a_10_n530# a1 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X102 full_adder_0/a_10_40# a1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X103 full_adder_0/a_1260_n530# a1 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X104 full_adder_0/a_1260_n530# b1 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X105 full_adder_0/a_760_40# b1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X106 full_adder_0/a_1260_40# b1 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X107 full_adder_0/a_2010_n530# full_adder_0/a_2670_n140# full_adder_0/a_2510_40# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X108 cout mux_2to1_4/a_2510_640# mux_2to1_4/in1 gnd sky130_fd_pr__nfet_01v8 ad=0.315 pd=3.2 as=0.315 ps=3.2 w=0.45 l=0.15
X109 cout mux_2to1_4/sel mux_2to1_4/in2 gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.45 l=0.15
X110 mux_2to1_4/a_2510_640# mux_2to1_4/sel gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X111 cout mux_2to1_4/sel mux_2to1_4/in1 vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=3.2 as=0.4725 ps=4.1 w=0.45 l=0.15
X112 cout mux_2to1_4/a_2510_640# mux_2to1_4/in2 vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.45 l=0.15
X113 mux_2to1_4/a_2510_640# mux_2to1_4/sel vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X114 full_adder_1/a_760_n530# b0 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X115 full_adder_1/a_510_n530# a0 full_adder_1/a_760_n530# gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X116 full_adder_0/cin full_adder_1/a_510_n530# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X117 full_adder_1/a_10_40# b0 vdd vdd sky130_fd_pr__pfet_01v8 ad=1.89 pd=12.9 as=0 ps=0 w=1.8 l=0.15
X118 full_adder_1/a_1260_40# cin0 vdd vdd sky130_fd_pr__pfet_01v8 ad=2.52 pd=17.2 as=0 ps=0 w=1.8 l=0.15
X119 full_adder_1/a_2260_40# a0 vdd vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=0 ps=0 w=1.8 l=0.15
X120 full_adder_1/a_10_n530# b0 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.945 pd=7.5 as=0 ps=0 w=0.9 l=0.15
X121 full_adder_1/a_510_n530# cin0 full_adder_1/a_10_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X122 full_adder_0/cin full_adder_1/a_510_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X123 full_adder_1/a_510_n530# a0 full_adder_1/a_760_40# vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=1.26 ps=8.6 w=1.8 l=0.15
X124 s0 full_adder_1/a_2010_n530# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X125 full_adder_1/a_2010_n530# full_adder_1/a_2670_n140# full_adder_1/a_2510_n530# gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0.63 ps=5 w=0.9 l=0.15
X126 s0 full_adder_1/a_2010_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X127 full_adder_1/a_1260_40# a0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X128 full_adder_1/a_510_n530# cin0 full_adder_1/a_10_40# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X129 full_adder_1/a_1260_n530# cin0 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.26 pd=10 as=0 ps=0 w=0.9 l=0.15
X130 full_adder_1/a_2010_n530# full_adder_1/a_510_n530# full_adder_1/a_1260_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X131 full_adder_1/a_2510_40# b0 full_adder_1/a_2260_40# vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=0 ps=0 w=1.8 l=0.15
X132 full_adder_1/a_2010_n530# full_adder_1/a_510_n530# full_adder_1/a_1260_40# vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=0 ps=0 w=1.8 l=0.15
X133 full_adder_1/a_2260_n530# a0 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X134 full_adder_1/a_2510_n530# b0 full_adder_1/a_2260_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X135 full_adder_1/a_10_n530# a0 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X136 full_adder_1/a_10_40# a0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X137 full_adder_1/a_1260_n530# a0 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X138 full_adder_1/a_1260_n530# b0 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X139 full_adder_1/a_760_40# b0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X140 full_adder_1/a_1260_40# b0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X141 full_adder_1/a_2010_n530# full_adder_1/a_2670_n140# full_adder_1/a_2510_40# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X142 full_adder_2/a_760_n530# b2 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X143 full_adder_2/a_510_n530# a2 full_adder_2/a_760_n530# gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X144 full_adder_4/cin full_adder_2/a_510_n530# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X145 full_adder_2/a_10_40# b2 vdd vdd sky130_fd_pr__pfet_01v8 ad=1.89 pd=12.9 as=0 ps=0 w=1.8 l=0.15
X146 full_adder_2/a_1260_40# full_adder_2/cin vdd vdd sky130_fd_pr__pfet_01v8 ad=2.52 pd=17.2 as=0 ps=0 w=1.8 l=0.15
X147 full_adder_2/a_2260_40# a2 vdd vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=0 ps=0 w=1.8 l=0.15
X148 full_adder_2/a_10_n530# b2 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.945 pd=7.5 as=0 ps=0 w=0.9 l=0.15
X149 full_adder_2/a_510_n530# full_adder_2/cin full_adder_2/a_10_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X150 full_adder_4/cin full_adder_2/a_510_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X151 full_adder_2/a_510_n530# a2 full_adder_2/a_760_40# vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=1.26 ps=8.6 w=1.8 l=0.15
X152 s2 full_adder_2/a_2010_n530# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X153 full_adder_2/a_2010_n530# full_adder_2/a_2670_n140# full_adder_2/a_2510_n530# gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0.63 ps=5 w=0.9 l=0.15
X154 s2 full_adder_2/a_2010_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X155 full_adder_2/a_1260_40# a2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X156 full_adder_2/a_510_n530# full_adder_2/cin full_adder_2/a_10_40# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X157 full_adder_2/a_1260_n530# full_adder_2/cin gnd gnd sky130_fd_pr__nfet_01v8 ad=1.26 pd=10 as=0 ps=0 w=0.9 l=0.15
X158 full_adder_2/a_2010_n530# full_adder_2/a_510_n530# full_adder_2/a_1260_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X159 full_adder_2/a_2510_40# b2 full_adder_2/a_2260_40# vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=0 ps=0 w=1.8 l=0.15
X160 full_adder_2/a_2010_n530# full_adder_2/a_510_n530# full_adder_2/a_1260_40# vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=0 ps=0 w=1.8 l=0.15
X161 full_adder_2/a_2260_n530# a2 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X162 full_adder_2/a_2510_n530# b2 full_adder_2/a_2260_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X163 full_adder_2/a_10_n530# a2 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X164 full_adder_2/a_10_40# a2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X165 full_adder_2/a_1260_n530# a2 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X166 full_adder_2/a_1260_n530# b2 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X167 full_adder_2/a_760_40# b2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X168 full_adder_2/a_1260_40# b2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X169 full_adder_2/a_2010_n530# full_adder_2/a_2670_n140# full_adder_2/a_2510_40# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X170 full_adder_3/a_760_n530# b7 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X171 full_adder_3/a_510_n530# a7 full_adder_3/a_760_n530# gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X172 mux_2to1_4/in1 full_adder_3/a_510_n530# full_adder_3/vdd full_adder_3/vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=5.04 ps=35.1 w=0.9 l=0.15
X173 full_adder_3/a_10_40# b7 full_adder_3/vdd full_adder_3/vdd sky130_fd_pr__pfet_01v8 ad=1.89 pd=12.9 as=0 ps=0 w=1.8 l=0.15
X174 full_adder_3/a_1260_40# full_adder_3/cin full_adder_3/vdd full_adder_3/vdd sky130_fd_pr__pfet_01v8 ad=2.52 pd=17.2 as=0 ps=0 w=1.8 l=0.15
X175 full_adder_3/a_2260_40# a7 full_adder_3/vdd full_adder_3/vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=0 ps=0 w=1.8 l=0.15
X176 full_adder_3/a_10_n530# b7 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.945 pd=7.5 as=0 ps=0 w=0.9 l=0.15
X177 full_adder_3/a_510_n530# full_adder_3/cin full_adder_3/a_10_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X178 mux_2to1_4/in1 full_adder_3/a_510_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.45 l=0.15
X179 full_adder_3/a_510_n530# a7 full_adder_3/a_760_40# full_adder_3/vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=1.26 ps=8.6 w=1.8 l=0.15
X180 mux_2to1_3/in1 full_adder_3/a_2010_n530# full_adder_3/vdd full_adder_3/vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X181 full_adder_3/a_2010_n530# full_adder_3/a_2670_n140# full_adder_3/a_2510_n530# gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0.63 ps=5 w=0.9 l=0.15
X182 mux_2to1_3/in1 full_adder_3/a_2010_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.45 l=0.15
X183 full_adder_3/a_1260_40# a7 full_adder_3/vdd full_adder_3/vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X184 full_adder_3/a_510_n530# full_adder_3/cin full_adder_3/a_10_40# full_adder_3/vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X185 full_adder_3/a_1260_n530# full_adder_3/cin gnd gnd sky130_fd_pr__nfet_01v8 ad=1.26 pd=10 as=0 ps=0 w=0.9 l=0.15
X186 full_adder_3/a_2010_n530# full_adder_3/a_510_n530# full_adder_3/a_1260_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X187 full_adder_3/a_2510_40# b7 full_adder_3/a_2260_40# full_adder_3/vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=0 ps=0 w=1.8 l=0.15
X188 full_adder_3/a_2010_n530# full_adder_3/a_510_n530# full_adder_3/a_1260_40# full_adder_3/vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=0 ps=0 w=1.8 l=0.15
X189 full_adder_3/a_2260_n530# a7 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X190 full_adder_3/a_2510_n530# b7 full_adder_3/a_2260_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X191 full_adder_3/a_10_n530# a7 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X192 full_adder_3/a_10_40# a7 full_adder_3/vdd full_adder_3/vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X193 full_adder_3/a_1260_n530# a7 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X194 full_adder_3/a_1260_n530# b7 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X195 full_adder_3/a_760_40# b7 full_adder_3/vdd full_adder_3/vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X196 full_adder_3/a_1260_40# b7 full_adder_3/vdd full_adder_3/vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X197 full_adder_3/a_2010_n530# full_adder_3/a_2670_n140# full_adder_3/a_2510_40# full_adder_3/vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X198 full_adder_4/a_760_n530# b3 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X199 full_adder_4/a_510_n530# a3 full_adder_4/a_760_n530# gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X200 mux_2to1_4/sel full_adder_4/a_510_n530# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X201 full_adder_4/a_10_40# b3 vdd vdd sky130_fd_pr__pfet_01v8 ad=1.89 pd=12.9 as=0 ps=0 w=1.8 l=0.15
X202 full_adder_4/a_1260_40# full_adder_4/cin vdd vdd sky130_fd_pr__pfet_01v8 ad=2.52 pd=17.2 as=0 ps=0 w=1.8 l=0.15
X203 full_adder_4/a_2260_40# a3 vdd vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=0 ps=0 w=1.8 l=0.15
X204 full_adder_4/a_10_n530# b3 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.945 pd=7.5 as=0 ps=0 w=0.9 l=0.15
X205 full_adder_4/a_510_n530# full_adder_4/cin full_adder_4/a_10_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X206 mux_2to1_4/sel full_adder_4/a_510_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X207 full_adder_4/a_510_n530# a3 full_adder_4/a_760_40# vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=1.26 ps=8.6 w=1.8 l=0.15
X208 s3 full_adder_4/a_2010_n530# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X209 full_adder_4/a_2010_n530# full_adder_4/a_2670_n140# full_adder_4/a_2510_n530# gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0.63 ps=5 w=0.9 l=0.15
X210 s3 full_adder_4/a_2010_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X211 full_adder_4/a_1260_40# a3 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X212 full_adder_4/a_510_n530# full_adder_4/cin full_adder_4/a_10_40# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X213 full_adder_4/a_1260_n530# full_adder_4/cin gnd gnd sky130_fd_pr__nfet_01v8 ad=1.26 pd=10 as=0 ps=0 w=0.9 l=0.15
X214 full_adder_4/a_2010_n530# full_adder_4/a_510_n530# full_adder_4/a_1260_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X215 full_adder_4/a_2510_40# b3 full_adder_4/a_2260_40# vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=0 ps=0 w=1.8 l=0.15
X216 full_adder_4/a_2010_n530# full_adder_4/a_510_n530# full_adder_4/a_1260_40# vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=0 ps=0 w=1.8 l=0.15
X217 full_adder_4/a_2260_n530# a3 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X218 full_adder_4/a_2510_n530# b3 full_adder_4/a_2260_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X219 full_adder_4/a_10_n530# a3 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X220 full_adder_4/a_10_40# a3 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X221 full_adder_4/a_1260_n530# a3 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X222 full_adder_4/a_1260_n530# b3 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X223 full_adder_4/a_760_40# b3 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X224 full_adder_4/a_1260_40# b3 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X225 full_adder_4/a_2010_n530# full_adder_4/a_2670_n140# full_adder_4/a_2510_40# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X226 full_adder_5/a_760_n530# b4 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X227 full_adder_5/a_510_n530# a4 full_adder_5/a_760_n530# gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X228 full_adder_6/cin full_adder_5/a_510_n530# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X229 full_adder_5/a_10_40# b4 vdd vdd sky130_fd_pr__pfet_01v8 ad=1.89 pd=12.9 as=0 ps=0 w=1.8 l=0.15
X230 full_adder_5/a_1260_40# cin0 vdd vdd sky130_fd_pr__pfet_01v8 ad=2.52 pd=17.2 as=0 ps=0 w=1.8 l=0.15
X231 full_adder_5/a_2260_40# a4 vdd vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=0 ps=0 w=1.8 l=0.15
X232 full_adder_5/a_10_n530# b4 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.945 pd=7.5 as=0 ps=0 w=0.9 l=0.15
X233 full_adder_5/a_510_n530# cin0 full_adder_5/a_10_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X234 full_adder_6/cin full_adder_5/a_510_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X235 full_adder_5/a_510_n530# a4 full_adder_5/a_760_40# vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=1.26 ps=8.6 w=1.8 l=0.15
X236 mux_2to1_0/in1 full_adder_5/a_2010_n530# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.4725 pd=4.1 as=0 ps=0 w=0.9 l=0.15
X237 full_adder_5/a_2010_n530# full_adder_5/a_2670_n140# full_adder_5/a_2510_n530# gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0.63 ps=5 w=0.9 l=0.15
X238 mux_2to1_0/in1 full_adder_5/a_2010_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.315 pd=3.2 as=0 ps=0 w=0.45 l=0.15
X239 full_adder_5/a_1260_40# a4 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X240 full_adder_5/a_510_n530# cin0 full_adder_5/a_10_40# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X241 full_adder_5/a_1260_n530# cin0 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.26 pd=10 as=0 ps=0 w=0.9 l=0.15
X242 full_adder_5/a_2010_n530# full_adder_5/a_510_n530# full_adder_5/a_1260_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X243 full_adder_5/a_2510_40# b4 full_adder_5/a_2260_40# vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=0 ps=0 w=1.8 l=0.15
X244 full_adder_5/a_2010_n530# full_adder_5/a_510_n530# full_adder_5/a_1260_40# vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=0 ps=0 w=1.8 l=0.15
X245 full_adder_5/a_2260_n530# a4 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X246 full_adder_5/a_2510_n530# b4 full_adder_5/a_2260_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X247 full_adder_5/a_10_n530# a4 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X248 full_adder_5/a_10_40# a4 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X249 full_adder_5/a_1260_n530# a4 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X250 full_adder_5/a_1260_n530# b4 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X251 full_adder_5/a_760_40# b4 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X252 full_adder_5/a_1260_40# b4 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X253 full_adder_5/a_2010_n530# full_adder_5/a_2670_n140# full_adder_5/a_2510_40# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X254 full_adder_6/a_760_n530# b5 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X255 full_adder_6/a_510_n530# a5 full_adder_6/a_760_n530# gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X256 full_adder_7/cin full_adder_6/a_510_n530# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X257 full_adder_6/a_10_40# b5 vdd vdd sky130_fd_pr__pfet_01v8 ad=1.89 pd=12.9 as=0 ps=0 w=1.8 l=0.15
X258 full_adder_6/a_1260_40# full_adder_6/cin vdd vdd sky130_fd_pr__pfet_01v8 ad=2.52 pd=17.2 as=0 ps=0 w=1.8 l=0.15
X259 full_adder_6/a_2260_40# a5 vdd vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=0 ps=0 w=1.8 l=0.15
X260 full_adder_6/a_10_n530# b5 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.945 pd=7.5 as=0 ps=0 w=0.9 l=0.15
X261 full_adder_6/a_510_n530# full_adder_6/cin full_adder_6/a_10_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X262 full_adder_7/cin full_adder_6/a_510_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X263 full_adder_6/a_510_n530# a5 full_adder_6/a_760_40# vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=1.26 ps=8.6 w=1.8 l=0.15
X264 mux_2to1_1/in1 full_adder_6/a_2010_n530# vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X265 full_adder_6/a_2010_n530# full_adder_6/a_2670_n140# full_adder_6/a_2510_n530# gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0.63 ps=5 w=0.9 l=0.15
X266 mux_2to1_1/in1 full_adder_6/a_2010_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.45 l=0.15
X267 full_adder_6/a_1260_40# a5 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X268 full_adder_6/a_510_n530# full_adder_6/cin full_adder_6/a_10_40# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X269 full_adder_6/a_1260_n530# full_adder_6/cin gnd gnd sky130_fd_pr__nfet_01v8 ad=1.26 pd=10 as=0 ps=0 w=0.9 l=0.15
X270 full_adder_6/a_2010_n530# full_adder_6/a_510_n530# full_adder_6/a_1260_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X271 full_adder_6/a_2510_40# b5 full_adder_6/a_2260_40# vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=0 ps=0 w=1.8 l=0.15
X272 full_adder_6/a_2010_n530# full_adder_6/a_510_n530# full_adder_6/a_1260_40# vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=0 ps=0 w=1.8 l=0.15
X273 full_adder_6/a_2260_n530# a5 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X274 full_adder_6/a_2510_n530# b5 full_adder_6/a_2260_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X275 full_adder_6/a_10_n530# a5 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X276 full_adder_6/a_10_40# a5 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X277 full_adder_6/a_1260_n530# a5 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X278 full_adder_6/a_1260_n530# b5 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X279 full_adder_6/a_760_40# b5 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X280 full_adder_6/a_1260_40# b5 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X281 full_adder_6/a_2010_n530# full_adder_6/a_2670_n140# full_adder_6/a_2510_40# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X282 full_adder_7/a_760_n530# b6 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X283 full_adder_7/a_510_n530# a6 full_adder_7/a_760_n530# gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X284 full_adder_3/cin full_adder_7/a_510_n530# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X285 full_adder_7/a_10_40# b6 vdd vdd sky130_fd_pr__pfet_01v8 ad=1.89 pd=12.9 as=0 ps=0 w=1.8 l=0.15
X286 full_adder_7/a_1260_40# full_adder_7/cin vdd vdd sky130_fd_pr__pfet_01v8 ad=2.52 pd=17.2 as=0 ps=0 w=1.8 l=0.15
X287 full_adder_7/a_2260_40# a6 vdd vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=0 ps=0 w=1.8 l=0.15
X288 full_adder_7/a_10_n530# b6 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.945 pd=7.5 as=0 ps=0 w=0.9 l=0.15
X289 full_adder_7/a_510_n530# full_adder_7/cin full_adder_7/a_10_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X290 full_adder_3/cin full_adder_7/a_510_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X291 full_adder_7/a_510_n530# a6 full_adder_7/a_760_40# vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=1.26 ps=8.6 w=1.8 l=0.15
X292 mux_2to1_2/in1 full_adder_7/a_2010_n530# vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X293 full_adder_7/a_2010_n530# full_adder_7/a_2670_n140# full_adder_7/a_2510_n530# gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0.63 ps=5 w=0.9 l=0.15
X294 mux_2to1_2/in1 full_adder_7/a_2010_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.45 l=0.15
X295 full_adder_7/a_1260_40# a6 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X296 full_adder_7/a_510_n530# full_adder_7/cin full_adder_7/a_10_40# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X297 full_adder_7/a_1260_n530# full_adder_7/cin gnd gnd sky130_fd_pr__nfet_01v8 ad=1.26 pd=10 as=0 ps=0 w=0.9 l=0.15
X298 full_adder_7/a_2010_n530# full_adder_7/a_510_n530# full_adder_7/a_1260_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X299 full_adder_7/a_2510_40# b6 full_adder_7/a_2260_40# vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=0 ps=0 w=1.8 l=0.15
X300 full_adder_7/a_2010_n530# full_adder_7/a_510_n530# full_adder_7/a_1260_40# vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=0 ps=0 w=1.8 l=0.15
X301 full_adder_7/a_2260_n530# a6 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X302 full_adder_7/a_2510_n530# b6 full_adder_7/a_2260_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X303 full_adder_7/a_10_n530# a6 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X304 full_adder_7/a_10_40# a6 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X305 full_adder_7/a_1260_n530# a6 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X306 full_adder_7/a_1260_n530# b6 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X307 full_adder_7/a_760_40# b6 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X308 full_adder_7/a_1260_40# b6 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X309 full_adder_7/a_2010_n530# full_adder_7/a_2670_n140# full_adder_7/a_2510_40# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X310 full_adder_8/a_760_n530# b5 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X311 full_adder_8/a_510_n530# a5 full_adder_8/a_760_n530# gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X312 full_adder_8/cout full_adder_8/a_510_n530# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X313 full_adder_8/a_10_40# b5 vdd vdd sky130_fd_pr__pfet_01v8 ad=1.89 pd=12.9 as=0 ps=0 w=1.8 l=0.15
X314 full_adder_8/a_1260_40# full_adder_8/cin vdd vdd sky130_fd_pr__pfet_01v8 ad=2.52 pd=17.2 as=0 ps=0 w=1.8 l=0.15
X315 full_adder_8/a_2260_40# a5 vdd vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=0 ps=0 w=1.8 l=0.15
X316 full_adder_8/a_10_n530# b5 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.945 pd=7.5 as=0 ps=0 w=0.9 l=0.15
X317 full_adder_8/a_510_n530# full_adder_8/cin full_adder_8/a_10_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X318 full_adder_8/cout full_adder_8/a_510_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X319 full_adder_8/a_510_n530# a5 full_adder_8/a_760_40# vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=1.26 ps=8.6 w=1.8 l=0.15
X320 mux_2to1_1/in2 full_adder_8/a_2010_n530# vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X321 full_adder_8/a_2010_n530# full_adder_8/a_2670_n140# full_adder_8/a_2510_n530# gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0.63 ps=5 w=0.9 l=0.15
X322 mux_2to1_1/in2 full_adder_8/a_2010_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.45 l=0.15
X323 full_adder_8/a_1260_40# a5 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X324 full_adder_8/a_510_n530# full_adder_8/cin full_adder_8/a_10_40# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X325 full_adder_8/a_1260_n530# full_adder_8/cin gnd gnd sky130_fd_pr__nfet_01v8 ad=1.26 pd=10 as=0 ps=0 w=0.9 l=0.15
X326 full_adder_8/a_2010_n530# full_adder_8/a_510_n530# full_adder_8/a_1260_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X327 full_adder_8/a_2510_40# b5 full_adder_8/a_2260_40# vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=0 ps=0 w=1.8 l=0.15
X328 full_adder_8/a_2010_n530# full_adder_8/a_510_n530# full_adder_8/a_1260_40# vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=0 ps=0 w=1.8 l=0.15
X329 full_adder_8/a_2260_n530# a5 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X330 full_adder_8/a_2510_n530# b5 full_adder_8/a_2260_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X331 full_adder_8/a_10_n530# a5 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X332 full_adder_8/a_10_40# a5 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X333 full_adder_8/a_1260_n530# a5 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X334 full_adder_8/a_1260_n530# b5 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X335 full_adder_8/a_760_40# b5 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X336 full_adder_8/a_1260_40# b5 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X337 full_adder_8/a_2010_n530# full_adder_8/a_2670_n140# full_adder_8/a_2510_40# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X338 full_adder_9/a_760_n530# b4 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X339 full_adder_9/a_510_n530# a4 full_adder_9/a_760_n530# gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X340 full_adder_8/cin full_adder_9/a_510_n530# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X341 full_adder_9/a_10_40# b4 vdd vdd sky130_fd_pr__pfet_01v8 ad=1.89 pd=12.9 as=0 ps=0 w=1.8 l=0.15
X342 full_adder_9/a_1260_40# cin1 vdd vdd sky130_fd_pr__pfet_01v8 ad=2.52 pd=17.2 as=0 ps=0 w=1.8 l=0.15
X343 full_adder_9/a_2260_40# a4 vdd vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=0 ps=0 w=1.8 l=0.15
X344 full_adder_9/a_10_n530# b4 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.945 pd=7.5 as=0 ps=0 w=0.9 l=0.15
X345 full_adder_9/a_510_n530# cin1 full_adder_9/a_10_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X346 full_adder_8/cin full_adder_9/a_510_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X347 full_adder_9/a_510_n530# a4 full_adder_9/a_760_40# vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=1.26 ps=8.6 w=1.8 l=0.15
X348 mux_2to1_0/in2 full_adder_9/a_2010_n530# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.4725 pd=4.1 as=0 ps=0 w=0.9 l=0.15
X349 full_adder_9/a_2010_n530# full_adder_9/a_2670_n140# full_adder_9/a_2510_n530# gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0.63 ps=5 w=0.9 l=0.15
X350 mux_2to1_0/in2 full_adder_9/a_2010_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.315 pd=3.2 as=0 ps=0 w=0.45 l=0.15
X351 full_adder_9/a_1260_40# a4 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X352 full_adder_9/a_510_n530# cin1 full_adder_9/a_10_40# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X353 full_adder_9/a_1260_n530# cin1 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.26 pd=10 as=0 ps=0 w=0.9 l=0.15
X354 full_adder_9/a_2010_n530# full_adder_9/a_510_n530# full_adder_9/a_1260_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X355 full_adder_9/a_2510_40# b4 full_adder_9/a_2260_40# vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=0 ps=0 w=1.8 l=0.15
X356 full_adder_9/a_2010_n530# full_adder_9/a_510_n530# full_adder_9/a_1260_40# vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=0 ps=0 w=1.8 l=0.15
X357 full_adder_9/a_2260_n530# a4 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X358 full_adder_9/a_2510_n530# b4 full_adder_9/a_2260_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X359 full_adder_9/a_10_n530# a4 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X360 full_adder_9/a_10_40# a4 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X361 full_adder_9/a_1260_n530# a4 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X362 full_adder_9/a_1260_n530# b4 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X363 full_adder_9/a_760_40# b4 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X364 full_adder_9/a_1260_40# b4 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X365 full_adder_9/a_2010_n530# full_adder_9/a_2670_n140# full_adder_9/a_2510_40# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
C0 b7 a7 18.335081f
C1 s5 s4 6.048123f
C2 mux_2to1_1/in1 mux_2to1_0/in1 12.358854f
C3 vdd a0 2.120752f
C4 mux_2to1_4/in1 mux_2to1_3/in2 3.99486f
C5 full_adder_3/vdd a7 2.112745f
C6 b5 a5 9.163856f
C7 full_adder_11/cin vdd 2.637957f
C8 vdd cin1 2.204039f
C9 b6 vdd 4.46876f
C10 s2 s1 2.236617f
C11 full_adder_7/cin vdd 2.63571f
C12 a6 b6 13.742169f
C13 vdd b0 2.142174f
C14 b4 cin1 2.868984f
C15 b0 cin0 2.618872f
C16 full_adder_8/cin vdd 2.640225f
C17 vdd mux_2to1_4/sel 3.484781f
C18 b2 a3 4.969382f
C19 full_adder_3/vdd full_adder_3/cin 2.432217f
C20 b2 full_adder_2/cin 2.030279f
C21 vdd cin0 4.406462f
C22 a6 vdd 4.75076f
C23 b2 a2 7.128378f
C24 s0 b7 4.435678f
C25 vdd b3 2.226849f
C26 vdd b7 2.330315f
C27 b4 vdd 4.29245f
C28 s5 s6 4.743982f
C29 b4 cin0 2.447221f
C30 vdd b5 4.513793f
C31 b1 a2 2.803949f
C32 a6 b5 5.052954f
C33 mux_2to1_0/in1 mux_2to1_4/sel 6.573423f
C34 full_adder_3/vdd b7 2.143207f
C35 vdd a4 4.369477f
C36 mux_2to1_0/in1 b7 4.436236f
C37 b4 a4 5.393144f
C38 b1 full_adder_0/cin 2.030289f
C39 vdd a3 2.28775f
C40 s0 s1 4.402915f
C41 vdd full_adder_2/cin 2.587097f
C42 b1 a1 4.892767f
C43 vdd a2 2.409542f
C44 mux_2to1_4/in1 mux_2to1_4/in2 2.720548f
C45 a3 b3 9.364401f
C46 mux_2to1_2/in1 mux_2to1_3/in1 5.389065f
C47 full_adder_8/cout vdd 2.636117f
C48 b6 a7 9.492191f
C49 vdd full_adder_0/cin 2.587147f
C50 vdd full_adder_4/cin 2.58683f
C51 s7 s6 3.439144f
C52 b2 vdd 2.249297f
C53 full_adder_4/cin b3 2.030272f
C54 vdd a1 2.930957f
C55 vdd a7 2.398573f
C56 vdd a5 5.547875f
C57 a0 b0 2.630623f
C58 mux_2to1_2/in1 mux_2to1_1/in1 8.667815f
C59 full_adder_6/cin vdd 2.640274f
C60 b1 vdd 2.313813f
C61 mux_2to1_4/sel gnd 13.61193f
C62 full_adder_9/a_510_n530# gnd 2.425663f 
C63 b4 gnd 3.171059f 
C64 a4 gnd 3.87003f
C65 full_adder_8/a_510_n530# gnd 2.427248f 
C66 b5 gnd 3.142176f 
C67 a5 gnd 3.600412f 
C68 full_adder_7/a_510_n530# gnd 2.425647f 
C69 full_adder_6/a_510_n530# gnd 2.427248f 
C70 full_adder_5/a_510_n530# gnd 2.425663f 
C71 full_adder_4/a_510_n530# gnd 2.425004f 
C72 full_adder_3/a_510_n530# gnd 2.425026f 
C73 full_adder_3/vdd gnd 9.098238f 
C74 full_adder_2/a_510_n530# gnd 2.425629f 
C75 full_adder_1/a_510_n530# gnd 2.425625f 
C76 full_adder_0/a_510_n530# gnd 2.425629f 
C77 vdd gnd 0.104133p 
C78 mux_2to1_1/in1 gnd 2.001458f 
C79 full_adder_11/a_510_n530# gnd 2.425026f 
C80 b7 gnd 3.825875f 
C81 a7 gnd 3.887742f 
C82 full_adder_10/a_510_n530# gnd 2.425647f 
C83 a6 gnd 3.705621f 


.end
