magic
tech sky130A
timestamp 1720436417
<< nwell >>
rect -30 90 130 285
<< nmos >>
rect 45 -25 60 20
<< pmos >>
rect 45 110 60 200
<< ndiff >>
rect 10 10 45 20
rect 10 -15 15 10
rect 35 -15 45 10
rect 10 -25 45 -15
rect 60 10 95 20
rect 60 -15 70 10
rect 90 -15 95 10
rect 60 -25 95 -15
<< pdiff >>
rect 10 190 45 200
rect 10 120 15 190
rect 35 120 45 190
rect 10 110 45 120
rect 60 190 95 200
rect 60 120 70 190
rect 90 120 95 190
rect 60 110 95 120
<< ndiffc >>
rect 15 -15 35 10
rect 70 -15 90 10
<< pdiffc >>
rect 15 120 35 190
rect 70 120 90 190
<< psubdiff >>
rect 0 -60 105 -55
rect 0 -80 15 -60
rect 35 -80 70 -60
rect 90 -80 105 -60
rect 0 -85 105 -80
<< nsubdiff >>
rect -10 255 110 260
rect -10 235 15 255
rect 35 235 70 255
rect 90 235 110 255
rect -10 230 110 235
<< psubdiffcont >>
rect 15 -80 35 -60
rect 70 -80 90 -60
<< nsubdiffcont >>
rect 15 235 35 255
rect 70 235 90 255
<< poly >>
rect 45 200 60 215
rect 45 70 60 110
rect 10 65 60 70
rect 10 45 20 65
rect 40 45 60 65
rect 10 40 60 45
rect 45 20 60 40
rect 45 -40 60 -25
<< polycont >>
rect 20 45 40 65
<< locali >>
rect -10 255 110 260
rect -10 235 15 255
rect 35 235 70 255
rect 90 235 110 255
rect -10 230 110 235
rect 15 200 35 230
rect 10 190 40 200
rect 10 120 15 190
rect 35 120 40 190
rect 10 110 40 120
rect 65 190 95 200
rect 65 120 70 190
rect 90 120 95 190
rect 65 110 95 120
rect 70 70 95 110
rect 10 65 50 70
rect 10 45 20 65
rect 40 45 50 65
rect 10 40 50 45
rect 70 65 120 70
rect 70 45 90 65
rect 110 45 120 65
rect 70 40 120 45
rect 70 20 95 40
rect 10 10 40 20
rect 10 -15 15 10
rect 35 -15 40 10
rect 10 -25 40 -15
rect 65 10 95 20
rect 65 -15 70 10
rect 90 -15 95 10
rect 65 -25 95 -15
rect 15 -55 35 -25
rect 0 -60 105 -55
rect 0 -80 15 -60
rect 35 -80 70 -60
rect 90 -80 105 -60
rect 0 -85 105 -80
<< viali >>
rect 70 235 90 255
rect 20 45 40 65
rect 90 45 110 65
rect 70 -80 90 -60
<< metal1 >>
rect -110 460 220 490
rect 60 255 100 460
rect 60 235 70 255
rect 90 235 100 255
rect 60 230 100 235
rect -110 65 50 70
rect -110 45 20 65
rect 40 45 50 65
rect -110 40 50 45
rect 80 65 180 70
rect 80 45 90 65
rect 110 45 180 65
rect 80 40 180 45
rect 60 -60 100 -55
rect 60 -80 70 -60
rect 90 -80 100 -60
rect 60 -230 100 -80
rect -110 -260 220 -230
<< labels >>
rlabel metal1 155 40 165 70 1 inv_outb
rlabel metal1 -80 40 -70 70 1 inv_in
rlabel metal1 80 470 80 470 1 vdd
rlabel metal1 90 -250 90 -250 1 gnd
<< end >>
