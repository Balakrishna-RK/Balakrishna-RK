magic
tech sky130A
timestamp 1720464950
<< nwell >>
rect 1180 440 1685 630
<< nmos >>
rect 1240 320 1255 365
rect 1395 320 1410 365
rect 1610 320 1625 365
<< pmos >>
rect 1240 460 1255 550
rect 1395 460 1410 505
rect 1610 460 1625 505
<< ndiff >>
rect 1205 355 1240 365
rect 1205 330 1210 355
rect 1230 330 1240 355
rect 1205 320 1240 330
rect 1255 355 1290 365
rect 1255 330 1265 355
rect 1285 330 1290 355
rect 1255 320 1290 330
rect 1360 355 1395 365
rect 1360 330 1365 355
rect 1385 330 1395 355
rect 1360 320 1395 330
rect 1410 355 1445 365
rect 1410 330 1420 355
rect 1440 330 1445 355
rect 1410 320 1445 330
rect 1575 355 1610 365
rect 1575 330 1580 355
rect 1600 330 1610 355
rect 1575 320 1610 330
rect 1625 355 1660 365
rect 1625 330 1635 355
rect 1655 330 1660 355
rect 1625 320 1660 330
<< pdiff >>
rect 1205 540 1240 550
rect 1205 520 1210 540
rect 1230 520 1240 540
rect 1205 490 1240 520
rect 1205 470 1210 490
rect 1230 470 1240 490
rect 1205 460 1240 470
rect 1255 540 1290 550
rect 1255 520 1265 540
rect 1285 520 1290 540
rect 1255 490 1290 520
rect 1255 470 1265 490
rect 1285 470 1290 490
rect 1255 460 1290 470
rect 1360 495 1395 505
rect 1360 470 1365 495
rect 1385 470 1395 495
rect 1360 460 1395 470
rect 1410 495 1445 505
rect 1410 470 1420 495
rect 1440 470 1445 495
rect 1410 460 1445 470
rect 1575 495 1610 505
rect 1575 470 1580 495
rect 1600 470 1610 495
rect 1575 460 1610 470
rect 1625 495 1660 505
rect 1625 470 1635 495
rect 1655 470 1660 495
rect 1625 460 1660 470
<< ndiffc >>
rect 1210 330 1230 355
rect 1265 330 1285 355
rect 1365 330 1385 355
rect 1420 330 1440 355
rect 1580 330 1600 355
rect 1635 330 1655 355
<< pdiffc >>
rect 1210 520 1230 540
rect 1210 470 1230 490
rect 1265 520 1285 540
rect 1265 470 1285 490
rect 1365 470 1385 495
rect 1420 470 1440 495
rect 1580 470 1600 495
rect 1635 470 1655 495
<< psubdiff >>
rect 1200 225 1295 230
rect 1200 205 1215 225
rect 1235 205 1260 225
rect 1280 205 1295 225
rect 1200 200 1295 205
rect 1355 225 1450 230
rect 1355 205 1370 225
rect 1390 205 1415 225
rect 1435 205 1450 225
rect 1355 200 1450 205
rect 1570 225 1665 230
rect 1570 205 1585 225
rect 1605 205 1630 225
rect 1650 205 1665 225
rect 1570 200 1665 205
<< nsubdiff >>
rect 1200 605 1295 610
rect 1200 585 1215 605
rect 1235 585 1260 605
rect 1280 585 1295 605
rect 1200 580 1295 585
rect 1355 605 1450 610
rect 1355 585 1370 605
rect 1390 585 1415 605
rect 1435 585 1450 605
rect 1355 580 1450 585
rect 1570 605 1665 610
rect 1570 585 1585 605
rect 1605 585 1630 605
rect 1650 585 1665 605
rect 1570 580 1665 585
<< psubdiffcont >>
rect 1215 205 1235 225
rect 1260 205 1280 225
rect 1370 205 1390 225
rect 1415 205 1435 225
rect 1585 205 1605 225
rect 1630 205 1650 225
<< nsubdiffcont >>
rect 1215 585 1235 605
rect 1260 585 1280 605
rect 1370 585 1390 605
rect 1415 585 1435 605
rect 1585 585 1605 605
rect 1630 585 1650 605
<< poly >>
rect 1240 550 1255 565
rect 1380 550 1420 555
rect 1380 530 1390 550
rect 1410 530 1420 550
rect 1380 525 1420 530
rect 1600 550 1640 555
rect 1600 530 1610 550
rect 1630 530 1640 550
rect 1600 525 1640 530
rect 1395 505 1410 525
rect 1610 505 1625 525
rect 1240 420 1255 460
rect 1395 445 1410 460
rect 1610 445 1625 460
rect 1205 415 1255 420
rect 1205 395 1215 415
rect 1235 395 1255 415
rect 1205 390 1255 395
rect 1240 365 1255 390
rect 1595 410 1635 415
rect 1595 390 1605 410
rect 1625 390 1635 410
rect 1595 385 1635 390
rect 1395 365 1410 380
rect 1610 365 1625 385
rect 1240 305 1255 320
rect 1395 300 1410 320
rect 1610 305 1625 320
rect 1385 295 1425 300
rect 1385 275 1395 295
rect 1415 275 1425 295
rect 1385 270 1425 275
<< polycont >>
rect 1390 530 1410 550
rect 1610 530 1630 550
rect 1215 395 1235 415
rect 1605 390 1625 410
rect 1395 275 1415 295
<< locali >>
rect 1560 700 1600 705
rect 1560 680 1570 700
rect 1590 680 1600 700
rect 1560 675 1600 680
rect 1570 655 1590 675
rect 1515 635 1590 655
rect 1200 605 1295 610
rect 1200 585 1215 605
rect 1235 585 1260 605
rect 1280 585 1295 605
rect 1200 580 1295 585
rect 1355 605 1450 610
rect 1355 585 1370 605
rect 1390 585 1415 605
rect 1435 585 1450 605
rect 1355 580 1450 585
rect 1210 550 1230 580
rect 1380 550 1420 555
rect 1205 540 1235 550
rect 1205 520 1210 540
rect 1230 520 1235 540
rect 1205 490 1235 520
rect 1205 470 1210 490
rect 1230 470 1235 490
rect 1205 460 1235 470
rect 1260 540 1290 550
rect 1260 520 1265 540
rect 1285 520 1290 540
rect 1380 530 1390 550
rect 1410 530 1420 550
rect 1380 525 1420 530
rect 1260 490 1290 520
rect 1260 470 1265 490
rect 1285 470 1290 490
rect 1260 460 1290 470
rect 1340 495 1390 505
rect 1340 470 1365 495
rect 1385 470 1390 495
rect 1340 460 1390 470
rect 1415 495 1465 505
rect 1415 470 1420 495
rect 1440 470 1465 495
rect 1415 460 1465 470
rect 1205 415 1245 420
rect 1205 395 1215 415
rect 1235 395 1245 415
rect 1205 390 1245 395
rect 1265 365 1285 460
rect 1340 420 1360 460
rect 1320 415 1360 420
rect 1320 395 1330 415
rect 1350 395 1360 415
rect 1320 390 1360 395
rect 1340 365 1360 390
rect 1445 365 1465 460
rect 1515 405 1535 635
rect 1570 605 1665 610
rect 1570 585 1585 605
rect 1605 585 1630 605
rect 1650 585 1665 605
rect 1570 580 1665 585
rect 1600 550 1640 555
rect 1600 530 1610 550
rect 1630 530 1640 550
rect 1600 525 1640 530
rect 1555 495 1605 505
rect 1555 470 1580 495
rect 1600 470 1605 495
rect 1555 460 1605 470
rect 1630 495 1680 505
rect 1630 470 1635 495
rect 1655 470 1680 495
rect 1630 460 1680 470
rect 1555 405 1575 460
rect 1515 385 1575 405
rect 1595 410 1635 415
rect 1595 390 1605 410
rect 1625 390 1635 410
rect 1595 385 1635 390
rect 1660 410 1680 460
rect 1740 410 1780 415
rect 1660 390 1750 410
rect 1770 390 1780 410
rect 1205 355 1235 365
rect 1205 330 1210 355
rect 1230 330 1235 355
rect 1205 320 1235 330
rect 1260 355 1290 365
rect 1260 330 1265 355
rect 1285 330 1290 355
rect 1260 320 1290 330
rect 1340 355 1390 365
rect 1340 330 1365 355
rect 1385 330 1390 355
rect 1340 320 1390 330
rect 1415 355 1465 365
rect 1415 330 1420 355
rect 1440 330 1465 355
rect 1415 320 1465 330
rect 1555 365 1575 385
rect 1660 365 1680 390
rect 1740 385 1780 390
rect 1555 355 1605 365
rect 1555 330 1580 355
rect 1600 330 1605 355
rect 1555 320 1605 330
rect 1630 355 1680 365
rect 1630 330 1635 355
rect 1655 330 1680 355
rect 1630 320 1680 330
rect 1210 230 1230 320
rect 1265 300 1285 320
rect 1255 295 1295 300
rect 1255 275 1265 295
rect 1285 275 1295 295
rect 1255 270 1295 275
rect 1385 295 1425 300
rect 1385 275 1395 295
rect 1415 275 1425 295
rect 1445 295 1465 320
rect 1660 295 1680 320
rect 1445 275 1680 295
rect 1385 270 1425 275
rect 1200 225 1295 230
rect 1200 205 1215 225
rect 1235 205 1260 225
rect 1280 205 1295 225
rect 1200 200 1295 205
rect 1355 225 1450 230
rect 1355 205 1370 225
rect 1390 205 1415 225
rect 1435 205 1450 225
rect 1355 200 1450 205
rect 1570 225 1665 230
rect 1570 205 1585 225
rect 1605 205 1630 225
rect 1650 205 1665 225
rect 1570 200 1665 205
<< viali >>
rect 1570 680 1590 700
rect 1260 585 1280 605
rect 1415 585 1435 605
rect 1390 530 1410 550
rect 1215 395 1235 415
rect 1330 395 1350 415
rect 1630 585 1650 605
rect 1610 530 1630 550
rect 1605 390 1625 410
rect 1750 390 1770 410
rect 1265 275 1285 295
rect 1395 275 1415 295
rect 1260 205 1280 225
rect 1415 205 1435 225
rect 1630 205 1650 225
<< metal1 >>
rect 1115 820 1650 840
rect 1155 700 1195 705
rect 1155 670 1160 700
rect 1190 670 1195 700
rect 1155 665 1195 670
rect 1165 415 1185 665
rect 1260 610 1280 820
rect 1300 750 1340 755
rect 1300 720 1305 750
rect 1335 720 1340 750
rect 1300 715 1340 720
rect 1250 605 1290 610
rect 1250 585 1260 605
rect 1280 585 1290 605
rect 1250 580 1290 585
rect 1310 420 1330 715
rect 1415 610 1435 820
rect 1560 800 1600 805
rect 1560 770 1565 800
rect 1595 770 1600 800
rect 1560 765 1600 770
rect 1570 705 1590 765
rect 1460 700 1500 705
rect 1460 670 1465 700
rect 1495 670 1500 700
rect 1560 700 1600 705
rect 1560 680 1570 700
rect 1590 680 1600 700
rect 1560 675 1600 680
rect 1460 665 1500 670
rect 1405 605 1445 610
rect 1405 585 1415 605
rect 1435 585 1445 605
rect 1405 580 1445 585
rect 1380 550 1420 555
rect 1470 550 1490 665
rect 1630 610 1650 820
rect 1620 605 1660 610
rect 1620 585 1630 605
rect 1650 585 1660 605
rect 1620 580 1660 585
rect 1600 550 1640 555
rect 1380 530 1390 550
rect 1410 530 1540 550
rect 1380 525 1420 530
rect 1205 415 1245 420
rect 1165 395 1215 415
rect 1235 395 1245 415
rect 1205 390 1245 395
rect 1310 415 1360 420
rect 1310 395 1330 415
rect 1350 395 1360 415
rect 1310 390 1360 395
rect 1520 405 1540 530
rect 1600 530 1610 550
rect 1630 530 1715 550
rect 1600 525 1640 530
rect 1595 410 1635 415
rect 1595 405 1605 410
rect 1520 390 1605 405
rect 1625 390 1635 410
rect 1520 385 1635 390
rect 1255 295 1295 300
rect 1385 295 1425 300
rect 1695 295 1715 530
rect 1740 410 1780 415
rect 1740 390 1750 410
rect 1770 390 1820 410
rect 1740 385 1780 390
rect 1255 275 1265 295
rect 1285 275 1395 295
rect 1415 275 1715 295
rect 1255 270 1295 275
rect 1385 270 1425 275
rect 1250 225 1290 230
rect 1250 205 1260 225
rect 1280 205 1290 225
rect 1250 200 1290 205
rect 1405 225 1445 230
rect 1405 205 1415 225
rect 1435 205 1445 225
rect 1405 200 1445 205
rect 1620 225 1660 230
rect 1620 205 1630 225
rect 1650 205 1660 225
rect 1620 200 1660 205
rect 1260 145 1280 200
rect 1415 145 1435 200
rect 1630 145 1650 200
rect 1115 125 1650 145
<< via1 >>
rect 1160 670 1190 700
rect 1305 720 1335 750
rect 1565 770 1595 800
rect 1465 670 1495 700
<< metal2 >>
rect 1560 800 1600 805
rect 1560 795 1565 800
rect 1115 775 1565 795
rect 1560 770 1565 775
rect 1595 770 1600 800
rect 1560 765 1600 770
rect 1300 750 1340 755
rect 1300 745 1305 750
rect 1115 725 1305 745
rect 1300 720 1305 725
rect 1335 720 1340 750
rect 1300 715 1340 720
rect 1155 700 1195 705
rect 1155 695 1160 700
rect 1115 675 1160 695
rect 1155 670 1160 675
rect 1190 695 1195 700
rect 1460 700 1500 705
rect 1460 695 1465 700
rect 1190 675 1465 695
rect 1190 670 1195 675
rect 1155 665 1195 670
rect 1460 670 1465 675
rect 1495 670 1500 700
rect 1460 665 1500 670
<< labels >>
rlabel metal2 1120 675 1130 695 1 sel
rlabel metal2 1120 725 1130 745 1 in1
rlabel metal2 1120 775 1130 795 1 in2
rlabel metal1 1320 130 1320 130 1 gnd
rlabel metal1 1240 830 1240 830 1 vdd
rlabel metal1 1800 390 1810 410 1 out
<< end >>
