* SPICE3 file created from mux_2to1.ext - technology: sky130A

Vin2 in2 GND PULSE(1.8 0 0 .1n .1n 10n 20n 8)
Vin1 in1 GND PULSE(1.8 0 0 .1n .1n 20n 40n 4)
Vsel sel GND PULSE(1.8 0 0 .1n .1n 20n 40n 2)
Vdd vdd GND 1.8

.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.tran .02ns 40ns
.save all


X0 out a_2510_640# in1 gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0.1575 ps=1.6 w=0.45 l=0.15
X1 out sel in2 gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0.1575 ps=1.6 w=0.45 l=0.15
X2 a_2510_640# sel gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0.1575 ps=1.6 w=0.45 l=0.15
X3 out sel in1 vdd sky130_fd_pr__pfet_01v8 ad=0.1575 pd=1.6 as=0.1575 ps=1.6 w=0.45 l=0.15
X4 out a_2510_640# in2 vdd sky130_fd_pr__pfet_01v8 ad=0.1575 pd=1.6 as=0.1575 ps=1.6 w=0.45 l=0.15
X5 a_2510_640# sel vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0.315 ps=2.5 w=0.9 l=0.15

.end
