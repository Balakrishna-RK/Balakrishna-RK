** sch_path: /home/krishna_rk/githubpro/cmoscharac/mos_charac/pmos/pmos_analysis.sch
**.subckt pmos_analysis
XM1 GND Vgs Vds Vds sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
Vgs Vds Vgs 0
Vds Vds GND 1.8
**** begin user architecture code

.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.dc Vds 0 1.8 0.1m Vgs 0 1.8 .3
.save all
.end

**** end user architecture code
**.ends
.GLOBAL GND
.end
