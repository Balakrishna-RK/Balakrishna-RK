* SPICE3 file created from carry_select_adder.ext - technology: sky130A

V17 cin0 GND 0
V18 cin1 GND 1.8
vdd vdd GND 1.8
V1 a0 GND PULSE(1.8 0 0 .1n .1n 80 90n 1)
V2 a1 GND PULSE(1.8 0 0 .1n .1n 40n 80n 2)
V3 a2 GND PULSE(1.8 0 0 .1n .1n 20n 40n 3)
V4 a3 GND PULSE(1.8 0 0 .1n .1n 10n 20n 4)
V5 a4 GND PULSE(0 1.8 0 .1n .1n 80 90n 1)
V6 a5 GND PULSE(0 1.8 0 .1n .1n 40n 80n 2)
V7 a6 GND PULSE(0 1.8 0 .1n .1n 20n 40n 3)
V8 a7 GND PULSE(0 1.8 0 .1n .1n 10n 20n 4)
V9 b0 GND PULSE(1.8 0 0 .1n .1n 80 90n 1)
V10 b1 GND PULSE(1.8 0 0 .1n .1n 40n 80n 2)
V11 b2 GND PULSE(1.8 0 0 .1n .1n 20n 40n 3)
V12 b3 GND PULSE(1.8 0 0 .1n .1n 10n 20n 4)
V13 b4 GND PULSE(0 1.8 0 .1n .1n 80 90n 1)
V14 b5 GND PULSE(0 1.8 0 .1n .1n 40n 80n 2)
V15 b6 GND PULSE(0 1.8 0 .1n .1n 20n 40n 3)
V16 b7 GND PULSE(0 1.8 0 .1n .1n 10n 20n 4)



.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.tran .02ns 80ns
.save all


X0 full_adder_10/a_3550_n440# full_adder_10/a_3010_n440# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0.315 ps=2.5 w=0.9 l=0.15
X1 full_adder_10/a_760_n530# b6 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.315 pd=2.5 as=0.315 ps=2.5 w=0.9 l=0.15
X2 full_adder_10/a_510_n530# a6 full_adder_10/a_760_n530# gnd sky130_fd_pr__nfet_01v8 ad=0.315 pd=2.5 as=0.315 ps=2.5 w=0.9 l=0.15
X3 full_adder_10/a_10_40# b6 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.63 pd=4.3 as=0.63 ps=4.3 w=1.8 l=0.15
X4 full_adder_10/a_3550_n440# full_adder_10/a_3010_n440# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0.1575 ps=1.6 w=0.45 l=0.15
X5 mux_2to1_2/in2 full_adder_10/a_3550_n440# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0.1575 ps=1.6 w=0.45 l=0.15
X6 full_adder_10/a_1260_40# full_adder_8/cout vdd vdd sky130_fd_pr__pfet_01v8 ad=0.63 pd=4.3 as=0.63 ps=4.3 w=1.8 l=0.15
X7 full_adder_10/a_2260_40# a6 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.945 pd=6.1 as=0.945 ps=6.1 w=2.7 l=0.15
X8 full_adder_10/a_10_n530# b6 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.315 pd=2.5 as=0.315 ps=2.5 w=0.9 l=0.15
X9 full_adder_10/a_510_n530# full_adder_8/cout full_adder_10/a_10_n530# gnd sky130_fd_pr__nfet_01v8 ad=0.315 pd=2.5 as=0.315 ps=2.5 w=0.9 l=0.15
X10 full_adder_10/a_510_n530# a6 full_adder_10/a_760_40# vdd sky130_fd_pr__pfet_01v8 ad=0.63 pd=4.3 as=0.63 ps=4.3 w=1.8 l=0.15
X11 full_adder_10/a_3010_n440# full_adder_10/a_2010_n530# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0.315 ps=2.5 w=0.9 l=0.15
X12 mux_2to1_2/in2 full_adder_10/a_3550_n440# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0.315 ps=2.5 w=0.9 l=0.15
X13 full_adder_11/cin full_adder_10/a_510_n530# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0.315 ps=2.5 w=0.9 l=0.15
X14 full_adder_10/a_2010_n530# full_adder_8/cout full_adder_10/a_2510_n620# gnd sky130_fd_pr__nfet_01v8 ad=0.4725 pd=3.4 as=0.4725 ps=3.4 w=1.35 l=0.15
X15 full_adder_10/a_3010_n440# full_adder_10/a_2010_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0.1575 ps=1.6 w=0.45 l=0.15
X16 full_adder_10/a_1260_40# a6 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.63 pd=4.3 as=0.63 ps=4.3 w=1.8 l=0.15
X17 full_adder_10/a_510_n530# full_adder_8/cout full_adder_10/a_10_40# vdd sky130_fd_pr__pfet_01v8 ad=0.63 pd=4.3 as=0.63 ps=4.3 w=1.8 l=0.15
X18 full_adder_10/a_1260_n530# full_adder_8/cout gnd gnd sky130_fd_pr__nfet_01v8 ad=0.315 pd=2.5 as=0.315 ps=2.5 w=0.9 l=0.15
X19 full_adder_10/a_2010_n530# full_adder_10/a_510_n530# full_adder_10/a_1260_n530# gnd sky130_fd_pr__nfet_01v8 ad=0.315 pd=2.5 as=0.315 ps=2.5 w=0.9 l=0.15
X20 full_adder_10/a_2510_40# b6 full_adder_10/a_2260_40# vdd sky130_fd_pr__pfet_01v8 ad=0.945 pd=6.1 as=0.945 ps=6.1 w=2.7 l=0.15
X21 full_adder_10/a_2010_n530# full_adder_10/a_510_n530# full_adder_10/a_1260_40# vdd sky130_fd_pr__pfet_01v8 ad=0.63 pd=4.3 as=0.63 ps=4.3 w=1.8 l=0.15
X22 full_adder_10/a_2260_n620# a6 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.4725 pd=3.4 as=0.4725 ps=3.4 w=1.35 l=0.15
X23 full_adder_10/a_2510_n620# b6 full_adder_10/a_2260_n620# gnd sky130_fd_pr__nfet_01v8 ad=0.4725 pd=3.4 as=0.4725 ps=3.4 w=1.35 l=0.15
X24 full_adder_11/cin full_adder_10/a_510_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0.1575 ps=1.6 w=0.45 l=0.15
X25 full_adder_10/a_10_n530# a6 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.315 pd=2.5 as=0.315 ps=2.5 w=0.9 l=0.15
X26 full_adder_10/a_10_40# a6 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.63 pd=4.3 as=0.63 ps=4.3 w=1.8 l=0.15
X27 full_adder_10/a_1260_n530# a6 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.315 pd=2.5 as=0.315 ps=2.5 w=0.9 l=0.15
X28 full_adder_10/a_1260_n530# b6 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.315 pd=2.5 as=0.315 ps=2.5 w=0.9 l=0.15
X29 full_adder_10/a_760_40# b6 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.63 pd=4.3 as=0.63 ps=4.3 w=1.8 l=0.15
X30 full_adder_10/a_1260_40# b6 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.63 pd=4.3 as=0.63 ps=4.3 w=1.8 l=0.15
X31 full_adder_10/a_2010_n530# full_adder_8/cout full_adder_10/a_2510_40# vdd sky130_fd_pr__pfet_01v8 ad=0.945 pd=6.1 as=0.945 ps=6.1 w=2.7 l=0.15
X32 full_adder_11/a_3550_n440# full_adder_11/a_3010_n440# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=76.23 ps=536.4 w=0.9 l=0.15
X33 full_adder_11/a_760_n530# b7 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=40.635 ps=338.6 w=0.9 l=0.15
X34 full_adder_11/a_510_n530# a7 full_adder_11/a_760_n530# gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X35 full_adder_11/a_10_40# b7 vdd vdd sky130_fd_pr__pfet_01v8 ad=1.89 pd=12.9 as=0 ps=0 w=1.8 l=0.15
X36 full_adder_11/a_3550_n440# full_adder_11/a_3010_n440# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X37 mux_2to1_3/in2 full_adder_11/a_3550_n440# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X38 full_adder_11/a_1260_40# full_adder_11/cin vdd vdd sky130_fd_pr__pfet_01v8 ad=2.52 pd=17.2 as=0 ps=0 w=1.8 l=0.15
X39 full_adder_11/a_2260_40# a7 vdd vdd sky130_fd_pr__pfet_01v8 ad=1.89 pd=12.2 as=0 ps=0 w=2.7 l=0.15
X40 full_adder_11/a_10_n530# b7 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.945 pd=7.5 as=0 ps=0 w=0.9 l=0.15
X41 full_adder_11/a_510_n530# full_adder_11/cin full_adder_11/a_10_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X42 full_adder_11/a_510_n530# a7 full_adder_11/a_760_40# vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=1.26 ps=8.6 w=1.8 l=0.15
X43 full_adder_11/a_3010_n440# full_adder_11/a_2010_n530# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X44 mux_2to1_3/in2 full_adder_11/a_3550_n440# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X45 mux_2to1_4/in2 full_adder_11/a_510_n530# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X46 full_adder_11/a_2010_n530# full_adder_11/cin full_adder_11/a_2510_n620# gnd sky130_fd_pr__nfet_01v8 ad=0.7875 pd=5.9 as=0.945 ps=6.8 w=1.35 l=0.15
X47 full_adder_11/a_3010_n440# full_adder_11/a_2010_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X48 full_adder_11/a_1260_40# a7 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X49 full_adder_11/a_510_n530# full_adder_11/cin full_adder_11/a_10_40# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X50 full_adder_11/a_1260_n530# full_adder_11/cin gnd gnd sky130_fd_pr__nfet_01v8 ad=1.26 pd=10 as=0 ps=0 w=0.9 l=0.15
X51 full_adder_11/a_2010_n530# full_adder_11/a_510_n530# full_adder_11/a_1260_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X52 full_adder_11/a_2510_40# b7 full_adder_11/a_2260_40# vdd sky130_fd_pr__pfet_01v8 ad=1.89 pd=12.2 as=0 ps=0 w=2.7 l=0.15
X53 full_adder_11/a_2010_n530# full_adder_11/a_510_n530# full_adder_11/a_1260_40# vdd sky130_fd_pr__pfet_01v8 ad=1.575 pd=10.4 as=0 ps=0 w=1.8 l=0.15
X54 full_adder_11/a_2260_n620# a7 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.945 pd=6.8 as=0 ps=0 w=1.35 l=0.15
X55 full_adder_11/a_2510_n620# b7 full_adder_11/a_2260_n620# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.35 l=0.15
X56 mux_2to1_4/in2 full_adder_11/a_510_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X57 full_adder_11/a_10_n530# a7 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X58 full_adder_11/a_10_40# a7 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X59 full_adder_11/a_1260_n530# a7 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X60 full_adder_11/a_1260_n530# b7 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X61 full_adder_11/a_760_40# b7 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X62 full_adder_11/a_1260_40# b7 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X63 full_adder_11/a_2010_n530# full_adder_11/cin full_adder_11/a_2510_40# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2.7 l=0.15
X64 mux_2to1_0/a_2720_340# mux_2to1_0/a_2510_640# mux_2to1_0/a_2820_860# vdd sky130_fd_pr__pfet_01v8 ad=0.63 pd=4.3 as=0.63 ps=4.3 w=1.8 l=0.15
X65 mux_2to1_0/a_2820_340# mux_2to1_4/sel mux_2to1_0/a_2720_340# gnd sky130_fd_pr__nfet_01v8 ad=0.315 pd=2.5 as=0.315 ps=2.5 w=0.9 l=0.15
X66 s4 mux_2to1_0/a_2720_340# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0.315 ps=2.5 w=0.9 l=0.15
X67 gnd mux_2to1_0/in2 mux_2to1_0/a_2820_340# gnd sky130_fd_pr__nfet_01v8 ad=0.315 pd=2.5 as=0.315 ps=2.5 w=0.9 l=0.15
X68 mux_2to1_0/a_2510_640# mux_2to1_4/sel gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0.1575 ps=1.6 w=0.45 l=0.15
X69 mux_2to1_0/a_3320_340# mux_2to1_0/a_2510_640# mux_2to1_0/a_2720_340# gnd sky130_fd_pr__nfet_01v8 ad=0.315 pd=2.5 as=0.315 ps=2.5 w=0.9 l=0.15
X70 mux_2to1_0/a_2720_340# vdd mux_2to1_0/a_2820_860# vdd sky130_fd_pr__pfet_01v8 ad=0.63 pd=4.3 as=0.63 ps=4.3 w=1.8 l=0.15
X71 s4 mux_2to1_0/a_2720_340# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0.1575 ps=1.6 w=0.45 l=0.15
X72 gnd vdd mux_2to1_0/a_3320_340# gnd sky130_fd_pr__nfet_01v8 ad=0.315 pd=2.5 as=0.315 ps=2.5 w=0.9 l=0.15
X73 mux_2to1_0/a_2820_860# mux_2to1_4/sel vdd vdd sky130_fd_pr__pfet_01v8 ad=0.63 pd=4.3 as=0.63 ps=4.3 w=1.8 l=0.15
X74 mux_2to1_0/a_2510_640# mux_2to1_4/sel vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0.315 ps=2.5 w=0.9 l=0.15
X75 mux_2to1_0/a_2820_860# mux_2to1_0/in2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0.63 pd=4.3 as=0.63 ps=4.3 w=1.8 l=0.15
X76 mux_2to1_1/a_2720_340# mux_2to1_1/a_2510_640# mux_2to1_1/a_2820_860# vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=2.52 ps=17.2 w=1.8 l=0.15
X77 mux_2to1_1/a_2820_340# mux_2to1_4/sel mux_2to1_1/a_2720_340# gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0.63 ps=5 w=0.9 l=0.15
X78 out mux_2to1_1/a_2720_340# vdd vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=10 as=0 ps=0 w=0.9 l=0.15
X79 gnd mux_2to1_1/in2 mux_2to1_1/a_2820_340# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X80 mux_2to1_1/a_2510_640# mux_2to1_4/sel gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X81 mux_2to1_1/a_3320_340# mux_2to1_1/a_2510_640# mux_2to1_1/a_2720_340# gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X82 mux_2to1_1/a_2720_340# vdd mux_2to1_1/a_2820_860# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X83 out mux_2to1_1/a_2720_340# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=6.4 as=0 ps=0 w=0.45 l=0.15
X84 gnd vdd mux_2to1_1/a_3320_340# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X85 mux_2to1_1/a_2820_860# mux_2to1_4/sel vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X86 mux_2to1_1/a_2510_640# mux_2to1_4/sel vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X87 mux_2to1_1/a_2820_860# mux_2to1_1/in2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X88 mux_2to1_2/a_2720_340# mux_2to1_2/a_2510_640# mux_2to1_2/a_2820_860# vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=2.52 ps=17.2 w=1.8 l=0.15
X89 mux_2to1_2/a_2820_340# mux_2to1_4/sel mux_2to1_2/a_2720_340# gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0.63 ps=5 w=0.9 l=0.15
X90 out mux_2to1_2/a_2720_340# vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X91 gnd mux_2to1_2/in2 mux_2to1_2/a_2820_340# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X92 mux_2to1_2/a_2510_640# mux_2to1_4/sel gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X93 mux_2to1_2/a_3320_340# mux_2to1_2/a_2510_640# mux_2to1_2/a_2720_340# gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X94 mux_2to1_2/a_2720_340# vdd mux_2to1_2/a_2820_860# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X95 out mux_2to1_2/a_2720_340# gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.45 l=0.15
X96 gnd vdd mux_2to1_2/a_3320_340# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X97 mux_2to1_2/a_2820_860# mux_2to1_4/sel vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X98 mux_2to1_2/a_2510_640# mux_2to1_4/sel vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X99 mux_2to1_2/a_2820_860# mux_2to1_2/in2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X100 full_adder_0/a_3550_n440# full_adder_0/a_3010_n440# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X101 full_adder_0/a_760_n530# full_adder_0/b gnd gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X102 full_adder_0/a_510_n530# full_adder_0/a full_adder_0/a_760_n530# gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X103 full_adder_0/a_10_40# full_adder_0/b vdd vdd sky130_fd_pr__pfet_01v8 ad=1.89 pd=12.9 as=0 ps=0 w=1.8 l=0.15
X104 full_adder_0/a_3550_n440# full_adder_0/a_3010_n440# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X105 s1 full_adder_0/a_3550_n440# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X106 full_adder_0/a_1260_40# full_adder_0/cin vdd vdd sky130_fd_pr__pfet_01v8 ad=2.52 pd=17.2 as=0 ps=0 w=1.8 l=0.15
X107 full_adder_0/a_2260_40# full_adder_0/a vdd vdd sky130_fd_pr__pfet_01v8 ad=1.89 pd=12.2 as=0 ps=0 w=2.7 l=0.15
X108 full_adder_0/a_10_n530# full_adder_0/b gnd gnd sky130_fd_pr__nfet_01v8 ad=0.945 pd=7.5 as=0 ps=0 w=0.9 l=0.15
X109 full_adder_0/a_510_n530# full_adder_0/cin full_adder_0/a_10_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X110 full_adder_0/a_510_n530# full_adder_0/a full_adder_0/a_760_40# vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=1.26 ps=8.6 w=1.8 l=0.15
X111 full_adder_0/a_3010_n440# full_adder_0/a_2010_n530# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X112 s1 full_adder_0/a_3550_n440# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X113 full_adder_2/cin full_adder_0/a_510_n530# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X114 full_adder_0/a_2010_n530# full_adder_0/cin full_adder_0/a_2510_n620# gnd sky130_fd_pr__nfet_01v8 ad=0.7875 pd=5.9 as=0.945 ps=6.8 w=1.35 l=0.15
X115 full_adder_0/a_3010_n440# full_adder_0/a_2010_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X116 full_adder_0/a_1260_40# full_adder_0/a vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X117 full_adder_0/a_510_n530# full_adder_0/cin full_adder_0/a_10_40# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X118 full_adder_0/a_1260_n530# full_adder_0/cin gnd gnd sky130_fd_pr__nfet_01v8 ad=1.26 pd=10 as=0 ps=0 w=0.9 l=0.15
X119 full_adder_0/a_2010_n530# full_adder_0/a_510_n530# full_adder_0/a_1260_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X120 full_adder_0/a_2510_40# full_adder_0/b full_adder_0/a_2260_40# vdd sky130_fd_pr__pfet_01v8 ad=1.89 pd=12.2 as=0 ps=0 w=2.7 l=0.15
X121 full_adder_0/a_2010_n530# full_adder_0/a_510_n530# full_adder_0/a_1260_40# vdd sky130_fd_pr__pfet_01v8 ad=1.575 pd=10.4 as=0 ps=0 w=1.8 l=0.15
X122 full_adder_0/a_2260_n620# full_adder_0/a gnd gnd sky130_fd_pr__nfet_01v8 ad=0.945 pd=6.8 as=0 ps=0 w=1.35 l=0.15
X123 full_adder_0/a_2510_n620# full_adder_0/b full_adder_0/a_2260_n620# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.35 l=0.15
X124 full_adder_2/cin full_adder_0/a_510_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X125 full_adder_0/a_10_n530# full_adder_0/a gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X126 full_adder_0/a_10_40# full_adder_0/a vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X127 full_adder_0/a_1260_n530# full_adder_0/a gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X128 full_adder_0/a_1260_n530# full_adder_0/b gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X129 full_adder_0/a_760_40# full_adder_0/b vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X130 full_adder_0/a_1260_40# full_adder_0/b vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X131 full_adder_0/a_2010_n530# full_adder_0/cin full_adder_0/a_2510_40# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2.7 l=0.15
X132 mux_2to1_3/a_2720_340# mux_2to1_3/a_2510_640# mux_2to1_3/a_2820_860# vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=2.52 ps=17.2 w=1.8 l=0.15
X133 mux_2to1_3/a_2820_340# mux_2to1_4/sel mux_2to1_3/a_2720_340# gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0.63 ps=5 w=0.9 l=0.15
X134 out mux_2to1_3/a_2720_340# vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X135 gnd mux_2to1_3/in2 mux_2to1_3/a_2820_340# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X136 mux_2to1_3/a_2510_640# mux_2to1_4/sel gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X137 mux_2to1_3/a_3320_340# mux_2to1_3/a_2510_640# mux_2to1_3/a_2720_340# gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X138 mux_2to1_3/a_2720_340# mux_2to1_3/in1 mux_2to1_3/a_2820_860# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X139 out mux_2to1_3/a_2720_340# gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.45 l=0.15
X140 gnd mux_2to1_3/in1 mux_2to1_3/a_3320_340# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X141 mux_2to1_3/a_2820_860# mux_2to1_4/sel vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X142 mux_2to1_3/a_2510_640# mux_2to1_4/sel vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X143 mux_2to1_3/a_2820_860# mux_2to1_3/in2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X144 mux_2to1_4/a_2720_340# mux_2to1_4/a_2510_640# mux_2to1_4/a_2820_860# vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=2.52 ps=17.2 w=1.8 l=0.15
X145 mux_2to1_4/a_2820_340# mux_2to1_4/sel mux_2to1_4/a_2720_340# gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0.63 ps=5 w=0.9 l=0.15
X146 out mux_2to1_4/a_2720_340# vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X147 gnd mux_2to1_4/in2 mux_2to1_4/a_2820_340# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X148 mux_2to1_4/a_2510_640# mux_2to1_4/sel gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X149 mux_2to1_4/a_3320_340# mux_2to1_4/a_2510_640# mux_2to1_4/a_2720_340# gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X150 mux_2to1_4/a_2720_340# mux_2to1_4/in1 mux_2to1_4/a_2820_860# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X151 out mux_2to1_4/a_2720_340# gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.45 l=0.15
X152 gnd mux_2to1_4/in1 mux_2to1_4/a_3320_340# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X153 mux_2to1_4/a_2820_860# mux_2to1_4/sel vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X154 mux_2to1_4/a_2510_640# mux_2to1_4/sel vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X155 mux_2to1_4/a_2820_860# mux_2to1_4/in2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X156 full_adder_1/a_3550_n440# full_adder_1/a_3010_n440# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X157 full_adder_1/a_760_n530# b0 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X158 full_adder_1/a_510_n530# a0 full_adder_1/a_760_n530# gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X159 full_adder_1/a_10_40# b0 vdd vdd sky130_fd_pr__pfet_01v8 ad=1.89 pd=12.9 as=0 ps=0 w=1.8 l=0.15
X160 full_adder_1/a_3550_n440# full_adder_1/a_3010_n440# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X161 s0 full_adder_1/a_3550_n440# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X162 full_adder_1/a_1260_40# cin0 vdd vdd sky130_fd_pr__pfet_01v8 ad=2.52 pd=17.2 as=0 ps=0 w=1.8 l=0.15
X163 full_adder_1/a_2260_40# a0 vdd vdd sky130_fd_pr__pfet_01v8 ad=1.89 pd=12.2 as=0 ps=0 w=2.7 l=0.15
X164 full_adder_1/a_10_n530# b0 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.945 pd=7.5 as=0 ps=0 w=0.9 l=0.15
X165 full_adder_1/a_510_n530# cin0 full_adder_1/a_10_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X166 full_adder_1/a_510_n530# a0 full_adder_1/a_760_40# vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=1.26 ps=8.6 w=1.8 l=0.15
X167 full_adder_1/a_3010_n440# full_adder_1/a_2010_n530# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X168 s0 full_adder_1/a_3550_n440# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X169 full_adder_0/cin full_adder_1/a_510_n530# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X170 full_adder_1/a_2010_n530# cin0 full_adder_1/a_2510_n620# gnd sky130_fd_pr__nfet_01v8 ad=0.7875 pd=5.9 as=0.945 ps=6.8 w=1.35 l=0.15
X171 full_adder_1/a_3010_n440# full_adder_1/a_2010_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X172 full_adder_1/a_1260_40# a0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X173 full_adder_1/a_510_n530# cin0 full_adder_1/a_10_40# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X174 full_adder_1/a_1260_n530# cin0 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.26 pd=10 as=0 ps=0 w=0.9 l=0.15
X175 full_adder_1/a_2010_n530# full_adder_1/a_510_n530# full_adder_1/a_1260_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X176 full_adder_1/a_2510_40# b0 full_adder_1/a_2260_40# vdd sky130_fd_pr__pfet_01v8 ad=1.89 pd=12.2 as=0 ps=0 w=2.7 l=0.15
X177 full_adder_1/a_2010_n530# full_adder_1/a_510_n530# full_adder_1/a_1260_40# vdd sky130_fd_pr__pfet_01v8 ad=1.575 pd=10.4 as=0 ps=0 w=1.8 l=0.15
X178 full_adder_1/a_2260_n620# a0 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.945 pd=6.8 as=0 ps=0 w=1.35 l=0.15
X179 full_adder_1/a_2510_n620# b0 full_adder_1/a_2260_n620# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.35 l=0.15
X180 full_adder_0/cin full_adder_1/a_510_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X181 full_adder_1/a_10_n530# a0 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X182 full_adder_1/a_10_40# a0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X183 full_adder_1/a_1260_n530# a0 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X184 full_adder_1/a_1260_n530# b0 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X185 full_adder_1/a_760_40# b0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X186 full_adder_1/a_1260_40# b0 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X187 full_adder_1/a_2010_n530# cin0 full_adder_1/a_2510_40# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2.7 l=0.15
X188 full_adder_3/a_3550_n440# full_adder_3/a_3010_n440# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X189 full_adder_3/a_760_n530# b7 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X190 full_adder_3/a_510_n530# a7 full_adder_3/a_760_n530# gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X191 full_adder_3/a_10_40# b7 vdd vdd sky130_fd_pr__pfet_01v8 ad=1.89 pd=12.9 as=0 ps=0 w=1.8 l=0.15
X192 full_adder_3/a_3550_n440# full_adder_3/a_3010_n440# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X193 mux_2to1_3/in1 full_adder_3/a_3550_n440# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X194 full_adder_3/a_1260_40# full_adder_3/cin vdd vdd sky130_fd_pr__pfet_01v8 ad=2.52 pd=17.2 as=0 ps=0 w=1.8 l=0.15
X195 full_adder_3/a_2260_40# a7 vdd vdd sky130_fd_pr__pfet_01v8 ad=1.89 pd=12.2 as=0 ps=0 w=2.7 l=0.15
X196 full_adder_3/a_10_n530# b7 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.945 pd=7.5 as=0 ps=0 w=0.9 l=0.15
X197 full_adder_3/a_510_n530# full_adder_3/cin full_adder_3/a_10_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X198 full_adder_3/a_510_n530# a7 full_adder_3/a_760_40# vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=1.26 ps=8.6 w=1.8 l=0.15
X199 full_adder_3/a_3010_n440# full_adder_3/a_2010_n530# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X200 mux_2to1_3/in1 full_adder_3/a_3550_n440# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X201 mux_2to1_4/in1 full_adder_3/a_510_n530# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X202 full_adder_3/a_2010_n530# full_adder_3/cin full_adder_3/a_2510_n620# gnd sky130_fd_pr__nfet_01v8 ad=0.7875 pd=5.9 as=0.945 ps=6.8 w=1.35 l=0.15
X203 full_adder_3/a_3010_n440# full_adder_3/a_2010_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X204 full_adder_3/a_1260_40# a7 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X205 full_adder_3/a_510_n530# full_adder_3/cin full_adder_3/a_10_40# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X206 full_adder_3/a_1260_n530# full_adder_3/cin gnd gnd sky130_fd_pr__nfet_01v8 ad=1.26 pd=10 as=0 ps=0 w=0.9 l=0.15
X207 full_adder_3/a_2010_n530# full_adder_3/a_510_n530# full_adder_3/a_1260_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X208 full_adder_3/a_2510_40# b7 full_adder_3/a_2260_40# vdd sky130_fd_pr__pfet_01v8 ad=1.89 pd=12.2 as=0 ps=0 w=2.7 l=0.15
X209 full_adder_3/a_2010_n530# full_adder_3/a_510_n530# full_adder_3/a_1260_40# vdd sky130_fd_pr__pfet_01v8 ad=1.575 pd=10.4 as=0 ps=0 w=1.8 l=0.15
X210 full_adder_3/a_2260_n620# a7 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.945 pd=6.8 as=0 ps=0 w=1.35 l=0.15
X211 full_adder_3/a_2510_n620# b7 full_adder_3/a_2260_n620# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.35 l=0.15
X212 mux_2to1_4/in1 full_adder_3/a_510_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X213 full_adder_3/a_10_n530# a7 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X214 full_adder_3/a_10_40# a7 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X215 full_adder_3/a_1260_n530# a7 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X216 full_adder_3/a_1260_n530# b7 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X217 full_adder_3/a_760_40# b7 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X218 full_adder_3/a_1260_40# b7 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X219 full_adder_3/a_2010_n530# full_adder_3/cin full_adder_3/a_2510_40# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2.7 l=0.15
X220 full_adder_2/a_3550_n440# full_adder_2/a_3010_n440# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X221 full_adder_2/a_760_n530# full_adder_2/b gnd gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X222 full_adder_2/a_510_n530# full_adder_2/a full_adder_2/a_760_n530# gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X223 full_adder_2/a_10_40# full_adder_2/b vdd vdd sky130_fd_pr__pfet_01v8 ad=1.89 pd=12.9 as=0 ps=0 w=1.8 l=0.15
X224 full_adder_2/a_3550_n440# full_adder_2/a_3010_n440# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X225 s2 full_adder_2/a_3550_n440# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X226 full_adder_2/a_1260_40# full_adder_2/cin vdd vdd sky130_fd_pr__pfet_01v8 ad=2.52 pd=17.2 as=0 ps=0 w=1.8 l=0.15
X227 full_adder_2/a_2260_40# full_adder_2/a vdd vdd sky130_fd_pr__pfet_01v8 ad=1.89 pd=12.2 as=0 ps=0 w=2.7 l=0.15
X228 full_adder_2/a_10_n530# full_adder_2/b gnd gnd sky130_fd_pr__nfet_01v8 ad=0.945 pd=7.5 as=0 ps=0 w=0.9 l=0.15
X229 full_adder_2/a_510_n530# full_adder_2/cin full_adder_2/a_10_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X230 full_adder_2/a_510_n530# full_adder_2/a full_adder_2/a_760_40# vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=1.26 ps=8.6 w=1.8 l=0.15
X231 full_adder_2/a_3010_n440# full_adder_2/a_2010_n530# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X232 s2 full_adder_2/a_3550_n440# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X233 full_adder_4/cin full_adder_2/a_510_n530# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X234 full_adder_2/a_2010_n530# full_adder_2/cin full_adder_2/a_2510_n620# gnd sky130_fd_pr__nfet_01v8 ad=0.7875 pd=5.9 as=0.945 ps=6.8 w=1.35 l=0.15
X235 full_adder_2/a_3010_n440# full_adder_2/a_2010_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X236 full_adder_2/a_1260_40# full_adder_2/a vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X237 full_adder_2/a_510_n530# full_adder_2/cin full_adder_2/a_10_40# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X238 full_adder_2/a_1260_n530# full_adder_2/cin gnd gnd sky130_fd_pr__nfet_01v8 ad=1.26 pd=10 as=0 ps=0 w=0.9 l=0.15
X239 full_adder_2/a_2010_n530# full_adder_2/a_510_n530# full_adder_2/a_1260_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X240 full_adder_2/a_2510_40# full_adder_2/b full_adder_2/a_2260_40# vdd sky130_fd_pr__pfet_01v8 ad=1.89 pd=12.2 as=0 ps=0 w=2.7 l=0.15
X241 full_adder_2/a_2010_n530# full_adder_2/a_510_n530# full_adder_2/a_1260_40# vdd sky130_fd_pr__pfet_01v8 ad=1.575 pd=10.4 as=0 ps=0 w=1.8 l=0.15
X242 full_adder_2/a_2260_n620# full_adder_2/a gnd gnd sky130_fd_pr__nfet_01v8 ad=0.945 pd=6.8 as=0 ps=0 w=1.35 l=0.15
X243 full_adder_2/a_2510_n620# full_adder_2/b full_adder_2/a_2260_n620# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.35 l=0.15
X244 full_adder_4/cin full_adder_2/a_510_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X245 full_adder_2/a_10_n530# full_adder_2/a gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X246 full_adder_2/a_10_40# full_adder_2/a vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X247 full_adder_2/a_1260_n530# full_adder_2/a gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X248 full_adder_2/a_1260_n530# full_adder_2/b gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X249 full_adder_2/a_760_40# full_adder_2/b vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X250 full_adder_2/a_1260_40# full_adder_2/b vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X251 full_adder_2/a_2010_n530# full_adder_2/cin full_adder_2/a_2510_40# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2.7 l=0.15
X252 full_adder_4/a_3550_n440# full_adder_4/a_3010_n440# full_adder_4/vdd full_adder_4/vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=5.985 ps=41.9 w=0.9 l=0.15
X253 full_adder_4/a_760_n530# b3 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X254 full_adder_4/a_510_n530# a3 full_adder_4/a_760_n530# gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X255 full_adder_4/a_10_40# b3 full_adder_4/vdd full_adder_4/vdd sky130_fd_pr__pfet_01v8 ad=1.89 pd=12.9 as=0 ps=0 w=1.8 l=0.15
X256 full_adder_4/a_3550_n440# full_adder_4/a_3010_n440# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X257 s3 full_adder_4/a_3550_n440# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X258 full_adder_4/a_1260_40# full_adder_4/cin full_adder_4/vdd full_adder_4/vdd sky130_fd_pr__pfet_01v8 ad=2.52 pd=17.2 as=0 ps=0 w=1.8 l=0.15
X259 full_adder_4/a_2260_40# a3 full_adder_4/vdd full_adder_4/vdd sky130_fd_pr__pfet_01v8 ad=1.89 pd=12.2 as=0 ps=0 w=2.7 l=0.15
X260 full_adder_4/a_10_n530# b3 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.945 pd=7.5 as=0 ps=0 w=0.9 l=0.15
X261 full_adder_4/a_510_n530# full_adder_4/cin full_adder_4/a_10_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X262 full_adder_4/a_510_n530# a3 full_adder_4/a_760_40# full_adder_4/vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=1.26 ps=8.6 w=1.8 l=0.15
X263 full_adder_4/a_3010_n440# full_adder_4/a_2010_n530# full_adder_4/vdd full_adder_4/vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X264 s3 full_adder_4/a_3550_n440# full_adder_4/vdd full_adder_4/vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X265 mux_2to1_4/sel full_adder_4/a_510_n530# full_adder_4/vdd full_adder_4/vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X266 full_adder_4/a_2010_n530# full_adder_4/cin full_adder_4/a_2510_n620# gnd sky130_fd_pr__nfet_01v8 ad=0.7875 pd=5.9 as=0.945 ps=6.8 w=1.35 l=0.15
X267 full_adder_4/a_3010_n440# full_adder_4/a_2010_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X268 full_adder_4/a_1260_40# a3 full_adder_4/vdd full_adder_4/vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X269 full_adder_4/a_510_n530# full_adder_4/cin full_adder_4/a_10_40# full_adder_4/vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X270 full_adder_4/a_1260_n530# full_adder_4/cin gnd gnd sky130_fd_pr__nfet_01v8 ad=1.26 pd=10 as=0 ps=0 w=0.9 l=0.15
X271 full_adder_4/a_2010_n530# full_adder_4/a_510_n530# full_adder_4/a_1260_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X272 full_adder_4/a_2510_40# b3 full_adder_4/a_2260_40# full_adder_4/vdd sky130_fd_pr__pfet_01v8 ad=1.89 pd=12.2 as=0 ps=0 w=2.7 l=0.15
X273 full_adder_4/a_2010_n530# full_adder_4/a_510_n530# full_adder_4/a_1260_40# full_adder_4/vdd sky130_fd_pr__pfet_01v8 ad=1.575 pd=10.4 as=0 ps=0 w=1.8 l=0.15
X274 full_adder_4/a_2260_n620# a3 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.945 pd=6.8 as=0 ps=0 w=1.35 l=0.15
X275 full_adder_4/a_2510_n620# b3 full_adder_4/a_2260_n620# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.35 l=0.15
X276 mux_2to1_4/sel full_adder_4/a_510_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X277 full_adder_4/a_10_n530# a3 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X278 full_adder_4/a_10_40# a3 full_adder_4/vdd full_adder_4/vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X279 full_adder_4/a_1260_n530# a3 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X280 full_adder_4/a_1260_n530# b3 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X281 full_adder_4/a_760_40# b3 full_adder_4/vdd full_adder_4/vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X282 full_adder_4/a_1260_40# b3 full_adder_4/vdd full_adder_4/vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X283 full_adder_4/a_2010_n530# full_adder_4/cin full_adder_4/a_2510_40# full_adder_4/vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2.7 l=0.15
X284 full_adder_5/a_3550_n440# full_adder_5/a_3010_n440# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X285 full_adder_5/a_760_n530# b4 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X286 full_adder_5/a_510_n530# a4 full_adder_5/a_760_n530# gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X287 full_adder_5/a_10_40# b4 vdd vdd sky130_fd_pr__pfet_01v8 ad=1.89 pd=12.9 as=0 ps=0 w=1.8 l=0.15
X288 full_adder_5/a_3550_n440# full_adder_5/a_3010_n440# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X289 vdd full_adder_5/a_3550_n440# gnd gnd sky130_fd_pr__nfet_01v8 ad=59.6225 pd=524.2 as=0 ps=0 w=0.45 l=0.15
X290 full_adder_5/a_1260_40# cin0 vdd vdd sky130_fd_pr__pfet_01v8 ad=2.52 pd=17.2 as=0 ps=0 w=1.8 l=0.15
X291 full_adder_5/a_2260_40# a4 vdd vdd sky130_fd_pr__pfet_01v8 ad=1.89 pd=12.2 as=0 ps=0 w=2.7 l=0.15
X292 full_adder_5/a_10_n530# b4 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.945 pd=7.5 as=0 ps=0 w=0.9 l=0.15
X293 full_adder_5/a_510_n530# cin0 full_adder_5/a_10_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X294 full_adder_5/a_510_n530# a4 full_adder_5/a_760_40# vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=1.26 ps=8.6 w=1.8 l=0.15
X295 full_adder_5/a_3010_n440# full_adder_5/a_2010_n530# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X296 vdd full_adder_5/a_3550_n440# vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X297 full_adder_6/cin full_adder_5/a_510_n530# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X298 full_adder_5/a_2010_n530# cin0 full_adder_5/a_2510_n620# gnd sky130_fd_pr__nfet_01v8 ad=0.7875 pd=5.9 as=0.945 ps=6.8 w=1.35 l=0.15
X299 full_adder_5/a_3010_n440# full_adder_5/a_2010_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X300 full_adder_5/a_1260_40# a4 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X301 full_adder_5/a_510_n530# cin0 full_adder_5/a_10_40# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X302 full_adder_5/a_1260_n530# cin0 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.26 pd=10 as=0 ps=0 w=0.9 l=0.15
X303 full_adder_5/a_2010_n530# full_adder_5/a_510_n530# full_adder_5/a_1260_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X304 full_adder_5/a_2510_40# b4 full_adder_5/a_2260_40# vdd sky130_fd_pr__pfet_01v8 ad=1.89 pd=12.2 as=0 ps=0 w=2.7 l=0.15
X305 full_adder_5/a_2010_n530# full_adder_5/a_510_n530# full_adder_5/a_1260_40# vdd sky130_fd_pr__pfet_01v8 ad=1.575 pd=10.4 as=0 ps=0 w=1.8 l=0.15
X306 full_adder_5/a_2260_n620# a4 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.945 pd=6.8 as=0 ps=0 w=1.35 l=0.15
X307 full_adder_5/a_2510_n620# b4 full_adder_5/a_2260_n620# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.35 l=0.15
X308 full_adder_6/cin full_adder_5/a_510_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X309 full_adder_5/a_10_n530# a4 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X310 full_adder_5/a_10_40# a4 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X311 full_adder_5/a_1260_n530# a4 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X312 full_adder_5/a_1260_n530# b4 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X313 full_adder_5/a_760_40# b4 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X314 full_adder_5/a_1260_40# b4 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X315 full_adder_5/a_2010_n530# cin0 full_adder_5/a_2510_40# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2.7 l=0.15
X316 full_adder_6/a_3550_n440# full_adder_6/a_3010_n440# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X317 full_adder_6/a_760_n530# b5 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X318 full_adder_6/a_510_n530# a5 full_adder_6/a_760_n530# gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X319 full_adder_6/a_10_40# b5 vdd vdd sky130_fd_pr__pfet_01v8 ad=1.89 pd=12.9 as=0 ps=0 w=1.8 l=0.15
X320 full_adder_6/a_3550_n440# full_adder_6/a_3010_n440# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X321 vdd full_adder_6/a_3550_n440# gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.45 l=0.15
X322 full_adder_6/a_1260_40# full_adder_6/cin vdd vdd sky130_fd_pr__pfet_01v8 ad=2.52 pd=17.2 as=0 ps=0 w=1.8 l=0.15
X323 full_adder_6/a_2260_40# a5 vdd vdd sky130_fd_pr__pfet_01v8 ad=1.89 pd=12.2 as=0 ps=0 w=2.7 l=0.15
X324 full_adder_6/a_10_n530# b5 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.945 pd=7.5 as=0 ps=0 w=0.9 l=0.15
X325 full_adder_6/a_510_n530# full_adder_6/cin full_adder_6/a_10_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X326 full_adder_6/a_510_n530# a5 full_adder_6/a_760_40# vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=1.26 ps=8.6 w=1.8 l=0.15
X327 full_adder_6/a_3010_n440# full_adder_6/a_2010_n530# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X328 vdd full_adder_6/a_3550_n440# vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X329 full_adder_7/cin full_adder_6/a_510_n530# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X330 full_adder_6/a_2010_n530# full_adder_6/cin full_adder_6/a_2510_n620# gnd sky130_fd_pr__nfet_01v8 ad=0.7875 pd=5.9 as=0.945 ps=6.8 w=1.35 l=0.15
X331 full_adder_6/a_3010_n440# full_adder_6/a_2010_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X332 full_adder_6/a_1260_40# a5 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X333 full_adder_6/a_510_n530# full_adder_6/cin full_adder_6/a_10_40# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X334 full_adder_6/a_1260_n530# full_adder_6/cin gnd gnd sky130_fd_pr__nfet_01v8 ad=1.26 pd=10 as=0 ps=0 w=0.9 l=0.15
X335 full_adder_6/a_2010_n530# full_adder_6/a_510_n530# full_adder_6/a_1260_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X336 full_adder_6/a_2510_40# b5 full_adder_6/a_2260_40# vdd sky130_fd_pr__pfet_01v8 ad=1.89 pd=12.2 as=0 ps=0 w=2.7 l=0.15
X337 full_adder_6/a_2010_n530# full_adder_6/a_510_n530# full_adder_6/a_1260_40# vdd sky130_fd_pr__pfet_01v8 ad=1.575 pd=10.4 as=0 ps=0 w=1.8 l=0.15
X338 full_adder_6/a_2260_n620# a5 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.945 pd=6.8 as=0 ps=0 w=1.35 l=0.15
X339 full_adder_6/a_2510_n620# b5 full_adder_6/a_2260_n620# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.35 l=0.15
X340 full_adder_7/cin full_adder_6/a_510_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X341 full_adder_6/a_10_n530# a5 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X342 full_adder_6/a_10_40# a5 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X343 full_adder_6/a_1260_n530# a5 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X344 full_adder_6/a_1260_n530# b5 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X345 full_adder_6/a_760_40# b5 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X346 full_adder_6/a_1260_40# b5 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X347 full_adder_6/a_2010_n530# full_adder_6/cin full_adder_6/a_2510_40# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2.7 l=0.15
X348 full_adder_7/a_3550_n440# full_adder_7/a_3010_n440# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X349 full_adder_7/a_760_n530# b6 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X350 full_adder_7/a_510_n530# a6 full_adder_7/a_760_n530# gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X351 full_adder_7/a_10_40# b6 vdd vdd sky130_fd_pr__pfet_01v8 ad=1.89 pd=12.9 as=0 ps=0 w=1.8 l=0.15
X352 full_adder_7/a_3550_n440# full_adder_7/a_3010_n440# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X353 vdd full_adder_7/a_3550_n440# gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.45 l=0.15
X354 full_adder_7/a_1260_40# full_adder_7/cin vdd vdd sky130_fd_pr__pfet_01v8 ad=2.52 pd=17.2 as=0 ps=0 w=1.8 l=0.15
X355 full_adder_7/a_2260_40# a6 vdd vdd sky130_fd_pr__pfet_01v8 ad=1.89 pd=12.2 as=0 ps=0 w=2.7 l=0.15
X356 full_adder_7/a_10_n530# b6 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.945 pd=7.5 as=0 ps=0 w=0.9 l=0.15
X357 full_adder_7/a_510_n530# full_adder_7/cin full_adder_7/a_10_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X358 full_adder_7/a_510_n530# a6 full_adder_7/a_760_40# vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=1.26 ps=8.6 w=1.8 l=0.15
X359 full_adder_7/a_3010_n440# full_adder_7/a_2010_n530# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X360 vdd full_adder_7/a_3550_n440# vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X361 full_adder_3/cin full_adder_7/a_510_n530# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X362 full_adder_7/a_2010_n530# full_adder_7/cin full_adder_7/a_2510_n620# gnd sky130_fd_pr__nfet_01v8 ad=0.7875 pd=5.9 as=0.945 ps=6.8 w=1.35 l=0.15
X363 full_adder_7/a_3010_n440# full_adder_7/a_2010_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X364 full_adder_7/a_1260_40# a6 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X365 full_adder_7/a_510_n530# full_adder_7/cin full_adder_7/a_10_40# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X366 full_adder_7/a_1260_n530# full_adder_7/cin gnd gnd sky130_fd_pr__nfet_01v8 ad=1.26 pd=10 as=0 ps=0 w=0.9 l=0.15
X367 full_adder_7/a_2010_n530# full_adder_7/a_510_n530# full_adder_7/a_1260_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X368 full_adder_7/a_2510_40# b6 full_adder_7/a_2260_40# vdd sky130_fd_pr__pfet_01v8 ad=1.89 pd=12.2 as=0 ps=0 w=2.7 l=0.15
X369 full_adder_7/a_2010_n530# full_adder_7/a_510_n530# full_adder_7/a_1260_40# vdd sky130_fd_pr__pfet_01v8 ad=1.575 pd=10.4 as=0 ps=0 w=1.8 l=0.15
X370 full_adder_7/a_2260_n620# a6 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.945 pd=6.8 as=0 ps=0 w=1.35 l=0.15
X371 full_adder_7/a_2510_n620# b6 full_adder_7/a_2260_n620# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.35 l=0.15
X372 full_adder_3/cin full_adder_7/a_510_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X373 full_adder_7/a_10_n530# a6 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X374 full_adder_7/a_10_40# a6 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X375 full_adder_7/a_1260_n530# a6 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X376 full_adder_7/a_1260_n530# b6 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X377 full_adder_7/a_760_40# b6 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X378 full_adder_7/a_1260_40# b6 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X379 full_adder_7/a_2010_n530# full_adder_7/cin full_adder_7/a_2510_40# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2.7 l=0.15
X380 full_adder_8/a_3550_n440# full_adder_8/a_3010_n440# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X381 full_adder_8/a_760_n530# b5 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X382 full_adder_8/a_510_n530# a5 full_adder_8/a_760_n530# gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X383 full_adder_8/a_10_40# b5 vdd vdd sky130_fd_pr__pfet_01v8 ad=1.89 pd=12.9 as=0 ps=0 w=1.8 l=0.15
X384 full_adder_8/a_3550_n440# full_adder_8/a_3010_n440# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X385 mux_2to1_1/in2 full_adder_8/a_3550_n440# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X386 full_adder_8/a_1260_40# full_adder_8/cin vdd vdd sky130_fd_pr__pfet_01v8 ad=2.52 pd=17.2 as=0 ps=0 w=1.8 l=0.15
X387 full_adder_8/a_2260_40# a5 vdd vdd sky130_fd_pr__pfet_01v8 ad=1.89 pd=12.2 as=0 ps=0 w=2.7 l=0.15
X388 full_adder_8/a_10_n530# b5 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.945 pd=7.5 as=0 ps=0 w=0.9 l=0.15
X389 full_adder_8/a_510_n530# full_adder_8/cin full_adder_8/a_10_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X390 full_adder_8/a_510_n530# a5 full_adder_8/a_760_40# vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=1.26 ps=8.6 w=1.8 l=0.15
X391 full_adder_8/a_3010_n440# full_adder_8/a_2010_n530# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X392 mux_2to1_1/in2 full_adder_8/a_3550_n440# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X393 full_adder_8/cout full_adder_8/a_510_n530# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X394 full_adder_8/a_2010_n530# full_adder_8/cin full_adder_8/a_2510_n620# gnd sky130_fd_pr__nfet_01v8 ad=0.7875 pd=5.9 as=0.945 ps=6.8 w=1.35 l=0.15
X395 full_adder_8/a_3010_n440# full_adder_8/a_2010_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X396 full_adder_8/a_1260_40# a5 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X397 full_adder_8/a_510_n530# full_adder_8/cin full_adder_8/a_10_40# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X398 full_adder_8/a_1260_n530# full_adder_8/cin gnd gnd sky130_fd_pr__nfet_01v8 ad=1.26 pd=10 as=0 ps=0 w=0.9 l=0.15
X399 full_adder_8/a_2010_n530# full_adder_8/a_510_n530# full_adder_8/a_1260_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X400 full_adder_8/a_2510_40# b5 full_adder_8/a_2260_40# vdd sky130_fd_pr__pfet_01v8 ad=1.89 pd=12.2 as=0 ps=0 w=2.7 l=0.15
X401 full_adder_8/a_2010_n530# full_adder_8/a_510_n530# full_adder_8/a_1260_40# vdd sky130_fd_pr__pfet_01v8 ad=1.575 pd=10.4 as=0 ps=0 w=1.8 l=0.15
X402 full_adder_8/a_2260_n620# a5 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.945 pd=6.8 as=0 ps=0 w=1.35 l=0.15
X403 full_adder_8/a_2510_n620# b5 full_adder_8/a_2260_n620# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.35 l=0.15
X404 full_adder_8/cout full_adder_8/a_510_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X405 full_adder_8/a_10_n530# a5 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X406 full_adder_8/a_10_40# a5 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X407 full_adder_8/a_1260_n530# a5 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X408 full_adder_8/a_1260_n530# b5 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X409 full_adder_8/a_760_40# b5 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X410 full_adder_8/a_1260_40# b5 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X411 full_adder_8/a_2010_n530# full_adder_8/cin full_adder_8/a_2510_40# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2.7 l=0.15
X412 full_adder_9/a_3550_n440# full_adder_9/a_3010_n440# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X413 full_adder_9/a_760_n530# b4 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X414 full_adder_9/a_510_n530# a4 full_adder_9/a_760_n530# gnd sky130_fd_pr__nfet_01v8 ad=0.63 pd=5 as=0 ps=0 w=0.9 l=0.15
X415 full_adder_9/a_10_40# b4 vdd vdd sky130_fd_pr__pfet_01v8 ad=1.89 pd=12.9 as=0 ps=0 w=1.8 l=0.15
X416 full_adder_9/a_3550_n440# full_adder_9/a_3010_n440# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X417 mux_2to1_0/in2 full_adder_9/a_3550_n440# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X418 full_adder_9/a_1260_40# cin1 vdd vdd sky130_fd_pr__pfet_01v8 ad=2.52 pd=17.2 as=0 ps=0 w=1.8 l=0.15
X419 full_adder_9/a_2260_40# a4 vdd vdd sky130_fd_pr__pfet_01v8 ad=1.89 pd=12.2 as=0 ps=0 w=2.7 l=0.15
X420 full_adder_9/a_10_n530# b4 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.945 pd=7.5 as=0 ps=0 w=0.9 l=0.15
X421 full_adder_9/a_510_n530# cin1 full_adder_9/a_10_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X422 full_adder_9/a_510_n530# a4 full_adder_9/a_760_40# vdd sky130_fd_pr__pfet_01v8 ad=1.26 pd=8.6 as=1.26 ps=8.6 w=1.8 l=0.15
X423 full_adder_9/a_3010_n440# full_adder_9/a_2010_n530# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X424 mux_2to1_0/in2 full_adder_9/a_3550_n440# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X425 full_adder_8/cin full_adder_9/a_510_n530# vdd vdd sky130_fd_pr__pfet_01v8 ad=0.315 pd=2.5 as=0 ps=0 w=0.9 l=0.15
X426 full_adder_9/a_2010_n530# cin1 full_adder_9/a_2510_n620# gnd sky130_fd_pr__nfet_01v8 ad=0.7875 pd=5.9 as=0.945 ps=6.8 w=1.35 l=0.15
X427 full_adder_9/a_3010_n440# full_adder_9/a_2010_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X428 full_adder_9/a_1260_40# a4 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X429 full_adder_9/a_510_n530# cin1 full_adder_9/a_10_40# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X430 full_adder_9/a_1260_n530# cin1 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.26 pd=10 as=0 ps=0 w=0.9 l=0.15
X431 full_adder_9/a_2010_n530# full_adder_9/a_510_n530# full_adder_9/a_1260_n530# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X432 full_adder_9/a_2510_40# b4 full_adder_9/a_2260_40# vdd sky130_fd_pr__pfet_01v8 ad=1.89 pd=12.2 as=0 ps=0 w=2.7 l=0.15
X433 full_adder_9/a_2010_n530# full_adder_9/a_510_n530# full_adder_9/a_1260_40# vdd sky130_fd_pr__pfet_01v8 ad=1.575 pd=10.4 as=0 ps=0 w=1.8 l=0.15
X434 full_adder_9/a_2260_n620# a4 gnd gnd sky130_fd_pr__nfet_01v8 ad=0.945 pd=6.8 as=0 ps=0 w=1.35 l=0.15
X435 full_adder_9/a_2510_n620# b4 full_adder_9/a_2260_n620# gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.35 l=0.15
X436 full_adder_8/cin full_adder_9/a_510_n530# gnd gnd sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.6 as=0 ps=0 w=0.45 l=0.15
X437 full_adder_9/a_10_n530# a4 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X438 full_adder_9/a_10_40# a4 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X439 full_adder_9/a_1260_n530# a4 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X440 full_adder_9/a_1260_n530# b4 gnd gnd sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.9 l=0.15
X441 full_adder_9/a_760_40# b4 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X442 full_adder_9/a_1260_40# b4 vdd vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=1.8 l=0.15
X443 full_adder_9/a_2010_n530# cin1 full_adder_9/a_2510_40# vdd sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=2.7 l=0.15
C0 full_adder_0/b full_adder_0/cin 2.175897f
C1 b5 full_adder_6/cin 2.175999f
C2 vdd full_adder_3/cin 3.110344f
C3 vdd a4 4.492331f
C4 b7 vdd 4.746863f
C5 vdd a7 5.032571f
C6 vdd full_adder_11/cin 2.988434f
C7 b3 full_adder_4/cin 2.175925f
C8 b3 full_adder_4/vdd 2.086557f
C9 b7 full_adder_3/cin 2.177865f
C10 vdd full_adder_0/cin 2.882514f
C11 b7 a7 20.622389f
C12 vdd full_adder_8/cout 2.995752f
C13 b7 full_adder_11/cin 2.17625f
C14 vdd full_adder_2/a 2.194557f
C15 vdd b6 4.526747f
C16 vdd a6 5.278062f
C17 full_adder_2/cin full_adder_2/b 2.175897f
C18 s1 s0 5.224577f
C19 b1 a2 3.05556f
C20 s1 s2 2.680423f
C21 a7 b6 10.770406f
C22 vdd full_adder_7/cin 3.113338f
C23 b5 full_adder_8/cin 2.174846f
C24 a1 b1 3.03111f
C25 a5 vdd 6.194f
C26 full_adder_8/cout b6 2.174836f
C27 mux_2to1_4/in2 mux_2to1_4/in1 2.497995f
C28 a3 full_adder_4/vdd 2.123355f
C29 a6 b6 15.273988f
C30 full_adder_2/b vdd 2.104858f
C31 vdd full_adder_6/cin 3.113338f
C32 mux_2to1_3/in1 mux_2to1_3/in2 4.545472f
C33 b2 a3 5.6f
C34 b5 vdd 4.532135f
C35 full_adder_7/cin b6 2.175999f
C36 b0 a0 2.670422f
C37 vdd a0 2.127173f
C38 b4 cin1 2.986482f
C39 full_adder_2/b full_adder_2/a 2.225328f
C40 a3 b3 10.508071f
C41 full_adder_0/b full_adder_0/a 2.225328f
C42 cin0 b4 2.564731f
C43 vdd cin1 2.452927f
C44 full_adder_8/cin vdd 2.997492f
C45 full_adder_2/cin vdd 2.882512f
C46 b5 a6 5.579248f
C47 cin0 b0 2.736369f
C48 cin0 vdd 4.89045f
C49 full_adder_0/b vdd 2.104858f
C50 vdd full_adder_0/a 2.194557f
C51 full_adder_4/vdd full_adder_4/cin 2.522835f
C52 b2 a2 5.64556f
C53 b4 vdd 4.190488f
C54 out s4 6.937213f
C55 vdd mux_2to1_2/in2 5.19392f
C56 out mux_2to1_4/sel 2.742471f
C57 s0 b7 5.146246f
C58 vdd mux_2to1_1/in2 5.469692f
C59 vdd b0 2.086375f
C60 b4 a4 5.472744f
C61 a5 b5 9.945868f
C62 vdd mux_2to1_0/in2 4.773131f
C63 vdd mux_2to1_4/sel 3.302925f
C64 full_adder_9/a_510_n530# gnd 2.263823f 
C65 b4 gnd 2.713483f 
C66 a4 gnd 3.403795f 
C67 full_adder_8/a_510_n530# gnd 2.263823f 
C68 b5 gnd 2.608924f 
C69 a5 gnd 3.201152f 
C70 full_adder_7/a_510_n530# gnd 2.263823f 
C71 full_adder_6/a_510_n530# gnd 2.263823f 
C72 full_adder_5/a_510_n530# gnd 2.263823f 
C73 full_adder_4/a_510_n530# gnd 2.2638f 
C74 full_adder_4/vdd gnd 13.145f 
C75 full_adder_4/cin gnd 2.069618f 
C76 full_adder_2/a_510_n530# gnd 2.2638f 
C77 full_adder_3/a_510_n530# gnd 2.263823f 
C78 full_adder_1/a_510_n530# gnd 2.2638f 
C79 mux_2to1_3/in1 gnd 2.484272f 
C80 full_adder_0/a_510_n530# gnd 2.2638f 
C81 out gnd 5.632544f 
C82 mux_2to1_4/sel gnd 13.906937f 
C83 vdd gnd 0.174676p 
C84 full_adder_11/a_510_n530# gnd 2.263823f
C85 b7 gnd 3.857558f 
C86 a7 gnd 3.677763f 
C87 full_adder_10/a_510_n530# gnd 2.263823f 
C88 b6 gnd 2.707542f 
C89 a6 gnd 3.372344f 

.end
