magic
tech sky130A
timestamp 1720949016
<< nwell >>
rect -70 -15 1960 475
rect 15 -20 230 -15
rect 1070 -20 1960 -15
<< nmos >>
rect -10 -265 5 -175
rect 115 -265 130 -175
rect 240 -265 255 -175
rect 365 -265 380 -175
rect 490 -265 505 -175
rect 615 -265 630 -175
rect 740 -265 755 -175
rect 865 -265 880 -175
rect 990 -265 1005 -175
rect 1115 -310 1130 -175
rect 1240 -310 1255 -175
rect 1365 -310 1380 -175
rect 1490 -220 1505 -175
rect 1630 -220 1645 -175
rect 1760 -220 1775 -175
rect 1885 -220 1900 -175
<< pmos >>
rect -10 20 5 200
rect 115 20 130 200
rect 240 20 255 200
rect 365 20 380 200
rect 490 20 505 200
rect 615 20 630 200
rect 740 20 755 200
rect 865 20 880 200
rect 990 20 1005 200
rect 1115 20 1130 290
rect 1240 20 1255 290
rect 1365 20 1380 290
rect 1490 20 1505 110
rect 1630 20 1645 110
rect 1760 20 1775 110
rect 1885 20 1900 110
<< ndiff >>
rect -45 -185 -10 -175
rect -45 -205 -40 -185
rect -20 -205 -10 -185
rect -45 -235 -10 -205
rect -45 -255 -40 -235
rect -20 -255 -10 -235
rect -45 -265 -10 -255
rect 5 -185 40 -175
rect 5 -205 15 -185
rect 35 -205 40 -185
rect 5 -235 40 -205
rect 5 -255 15 -235
rect 35 -255 40 -235
rect 5 -265 40 -255
rect 80 -185 115 -175
rect 80 -205 85 -185
rect 105 -205 115 -185
rect 80 -235 115 -205
rect 80 -255 85 -235
rect 105 -255 115 -235
rect 80 -265 115 -255
rect 130 -185 165 -175
rect 130 -205 140 -185
rect 160 -205 165 -185
rect 130 -235 165 -205
rect 130 -255 140 -235
rect 160 -255 165 -235
rect 130 -265 165 -255
rect 205 -185 240 -175
rect 205 -205 210 -185
rect 230 -205 240 -185
rect 205 -235 240 -205
rect 205 -255 210 -235
rect 230 -255 240 -235
rect 205 -265 240 -255
rect 255 -185 290 -175
rect 255 -205 265 -185
rect 285 -205 290 -185
rect 255 -235 290 -205
rect 255 -255 265 -235
rect 285 -255 290 -235
rect 255 -265 290 -255
rect 330 -185 365 -175
rect 330 -205 335 -185
rect 355 -205 365 -185
rect 330 -235 365 -205
rect 330 -255 335 -235
rect 355 -255 365 -235
rect 330 -265 365 -255
rect 380 -185 415 -175
rect 380 -205 390 -185
rect 410 -205 415 -185
rect 380 -235 415 -205
rect 380 -255 390 -235
rect 410 -255 415 -235
rect 380 -265 415 -255
rect 455 -185 490 -175
rect 455 -205 460 -185
rect 480 -205 490 -185
rect 455 -235 490 -205
rect 455 -255 460 -235
rect 480 -255 490 -235
rect 455 -265 490 -255
rect 505 -185 540 -175
rect 505 -205 515 -185
rect 535 -205 540 -185
rect 505 -235 540 -205
rect 505 -255 515 -235
rect 535 -255 540 -235
rect 505 -265 540 -255
rect 580 -185 615 -175
rect 580 -205 585 -185
rect 605 -205 615 -185
rect 580 -235 615 -205
rect 580 -255 585 -235
rect 605 -255 615 -235
rect 580 -265 615 -255
rect 630 -185 665 -175
rect 630 -205 640 -185
rect 660 -205 665 -185
rect 630 -235 665 -205
rect 630 -255 640 -235
rect 660 -255 665 -235
rect 630 -265 665 -255
rect 705 -185 740 -175
rect 705 -205 710 -185
rect 730 -205 740 -185
rect 705 -235 740 -205
rect 705 -255 710 -235
rect 730 -255 740 -235
rect 705 -265 740 -255
rect 755 -185 790 -175
rect 755 -205 765 -185
rect 785 -205 790 -185
rect 755 -235 790 -205
rect 755 -255 765 -235
rect 785 -255 790 -235
rect 755 -265 790 -255
rect 830 -185 865 -175
rect 830 -205 835 -185
rect 855 -205 865 -185
rect 830 -235 865 -205
rect 830 -255 835 -235
rect 855 -255 865 -235
rect 830 -265 865 -255
rect 880 -185 915 -175
rect 880 -205 890 -185
rect 910 -205 915 -185
rect 880 -235 915 -205
rect 880 -255 890 -235
rect 910 -255 915 -235
rect 880 -265 915 -255
rect 955 -185 990 -175
rect 955 -205 960 -185
rect 980 -205 990 -185
rect 955 -235 990 -205
rect 955 -255 960 -235
rect 980 -255 990 -235
rect 955 -265 990 -255
rect 1005 -185 1040 -175
rect 1005 -205 1015 -185
rect 1035 -205 1040 -185
rect 1005 -235 1040 -205
rect 1005 -255 1015 -235
rect 1035 -255 1040 -235
rect 1005 -265 1040 -255
rect 1080 -185 1115 -175
rect 1080 -205 1085 -185
rect 1105 -205 1115 -185
rect 1080 -235 1115 -205
rect 1080 -255 1085 -235
rect 1105 -255 1115 -235
rect 1080 -280 1115 -255
rect 1080 -300 1085 -280
rect 1105 -300 1115 -280
rect 1080 -310 1115 -300
rect 1130 -185 1165 -175
rect 1130 -205 1140 -185
rect 1160 -205 1165 -185
rect 1130 -235 1165 -205
rect 1130 -255 1140 -235
rect 1160 -255 1165 -235
rect 1130 -280 1165 -255
rect 1130 -300 1140 -280
rect 1160 -300 1165 -280
rect 1130 -310 1165 -300
rect 1205 -185 1240 -175
rect 1205 -205 1210 -185
rect 1230 -205 1240 -185
rect 1205 -235 1240 -205
rect 1205 -255 1210 -235
rect 1230 -255 1240 -235
rect 1205 -280 1240 -255
rect 1205 -300 1210 -280
rect 1230 -300 1240 -280
rect 1205 -310 1240 -300
rect 1255 -185 1290 -175
rect 1255 -205 1265 -185
rect 1285 -205 1290 -185
rect 1255 -235 1290 -205
rect 1255 -255 1265 -235
rect 1285 -255 1290 -235
rect 1255 -280 1290 -255
rect 1255 -300 1265 -280
rect 1285 -300 1290 -280
rect 1255 -310 1290 -300
rect 1330 -185 1365 -175
rect 1330 -205 1335 -185
rect 1355 -205 1365 -185
rect 1330 -235 1365 -205
rect 1330 -255 1335 -235
rect 1355 -255 1365 -235
rect 1330 -280 1365 -255
rect 1330 -300 1335 -280
rect 1355 -300 1365 -280
rect 1330 -310 1365 -300
rect 1380 -185 1415 -175
rect 1380 -205 1390 -185
rect 1410 -205 1415 -185
rect 1380 -235 1415 -205
rect 1455 -185 1490 -175
rect 1455 -210 1460 -185
rect 1480 -210 1490 -185
rect 1455 -220 1490 -210
rect 1505 -185 1540 -175
rect 1505 -210 1515 -185
rect 1535 -210 1540 -185
rect 1505 -220 1540 -210
rect 1595 -185 1630 -175
rect 1595 -210 1600 -185
rect 1620 -210 1630 -185
rect 1595 -220 1630 -210
rect 1645 -185 1680 -175
rect 1645 -210 1655 -185
rect 1675 -210 1680 -185
rect 1645 -220 1680 -210
rect 1725 -185 1760 -175
rect 1725 -210 1730 -185
rect 1750 -210 1760 -185
rect 1725 -220 1760 -210
rect 1775 -185 1810 -175
rect 1775 -210 1785 -185
rect 1805 -210 1810 -185
rect 1775 -220 1810 -210
rect 1850 -185 1885 -175
rect 1850 -210 1855 -185
rect 1875 -210 1885 -185
rect 1850 -220 1885 -210
rect 1900 -185 1935 -175
rect 1900 -210 1910 -185
rect 1930 -210 1935 -185
rect 1900 -220 1935 -210
rect 1380 -255 1390 -235
rect 1410 -255 1415 -235
rect 1380 -280 1415 -255
rect 1380 -300 1390 -280
rect 1410 -300 1415 -280
rect 1380 -310 1415 -300
<< pdiff >>
rect 1080 280 1115 290
rect 1080 260 1085 280
rect 1105 260 1115 280
rect 1080 240 1115 260
rect 1080 220 1085 240
rect 1105 220 1115 240
rect -45 190 -10 200
rect -45 170 -40 190
rect -20 170 -10 190
rect -45 140 -10 170
rect -45 120 -40 140
rect -20 120 -10 140
rect -45 100 -10 120
rect -45 80 -40 100
rect -20 80 -10 100
rect -45 50 -10 80
rect -45 30 -40 50
rect -20 30 -10 50
rect -45 20 -10 30
rect 5 190 40 200
rect 5 170 15 190
rect 35 170 40 190
rect 5 140 40 170
rect 5 120 15 140
rect 35 120 40 140
rect 5 100 40 120
rect 5 80 15 100
rect 35 80 40 100
rect 5 50 40 80
rect 5 30 15 50
rect 35 30 40 50
rect 5 20 40 30
rect 80 190 115 200
rect 80 170 85 190
rect 105 170 115 190
rect 80 140 115 170
rect 80 120 85 140
rect 105 120 115 140
rect 80 100 115 120
rect 80 80 85 100
rect 105 80 115 100
rect 80 50 115 80
rect 80 30 85 50
rect 105 30 115 50
rect 80 20 115 30
rect 130 190 165 200
rect 130 170 140 190
rect 160 170 165 190
rect 130 140 165 170
rect 130 120 140 140
rect 160 120 165 140
rect 130 100 165 120
rect 130 80 140 100
rect 160 80 165 100
rect 130 50 165 80
rect 130 30 140 50
rect 160 30 165 50
rect 130 20 165 30
rect 205 190 240 200
rect 205 170 210 190
rect 230 170 240 190
rect 205 140 240 170
rect 205 120 210 140
rect 230 120 240 140
rect 205 100 240 120
rect 205 80 210 100
rect 230 80 240 100
rect 205 50 240 80
rect 205 30 210 50
rect 230 30 240 50
rect 205 20 240 30
rect 255 190 290 200
rect 255 170 265 190
rect 285 170 290 190
rect 255 140 290 170
rect 255 120 265 140
rect 285 120 290 140
rect 255 100 290 120
rect 255 80 265 100
rect 285 80 290 100
rect 255 50 290 80
rect 255 30 265 50
rect 285 30 290 50
rect 255 20 290 30
rect 330 190 365 200
rect 330 170 335 190
rect 355 170 365 190
rect 330 140 365 170
rect 330 120 335 140
rect 355 120 365 140
rect 330 100 365 120
rect 330 80 335 100
rect 355 80 365 100
rect 330 50 365 80
rect 330 30 335 50
rect 355 30 365 50
rect 330 20 365 30
rect 380 190 415 200
rect 380 170 390 190
rect 410 170 415 190
rect 380 140 415 170
rect 380 120 390 140
rect 410 120 415 140
rect 380 100 415 120
rect 380 80 390 100
rect 410 80 415 100
rect 380 50 415 80
rect 380 30 390 50
rect 410 30 415 50
rect 380 20 415 30
rect 455 190 490 200
rect 455 170 460 190
rect 480 170 490 190
rect 455 140 490 170
rect 455 120 460 140
rect 480 120 490 140
rect 455 100 490 120
rect 455 80 460 100
rect 480 80 490 100
rect 455 50 490 80
rect 455 30 460 50
rect 480 30 490 50
rect 455 20 490 30
rect 505 190 540 200
rect 505 170 515 190
rect 535 170 540 190
rect 505 140 540 170
rect 505 120 515 140
rect 535 120 540 140
rect 505 100 540 120
rect 505 80 515 100
rect 535 80 540 100
rect 505 50 540 80
rect 505 30 515 50
rect 535 30 540 50
rect 505 20 540 30
rect 580 190 615 200
rect 580 170 585 190
rect 605 170 615 190
rect 580 140 615 170
rect 580 120 585 140
rect 605 120 615 140
rect 580 100 615 120
rect 580 80 585 100
rect 605 80 615 100
rect 580 50 615 80
rect 580 30 585 50
rect 605 30 615 50
rect 580 20 615 30
rect 630 190 665 200
rect 630 170 640 190
rect 660 170 665 190
rect 630 140 665 170
rect 630 120 640 140
rect 660 120 665 140
rect 630 100 665 120
rect 630 80 640 100
rect 660 80 665 100
rect 630 50 665 80
rect 630 30 640 50
rect 660 30 665 50
rect 630 20 665 30
rect 705 190 740 200
rect 705 170 710 190
rect 730 170 740 190
rect 705 140 740 170
rect 705 120 710 140
rect 730 120 740 140
rect 705 100 740 120
rect 705 80 710 100
rect 730 80 740 100
rect 705 50 740 80
rect 705 30 710 50
rect 730 30 740 50
rect 705 20 740 30
rect 755 190 790 200
rect 755 170 765 190
rect 785 170 790 190
rect 755 140 790 170
rect 755 120 765 140
rect 785 120 790 140
rect 755 100 790 120
rect 755 80 765 100
rect 785 80 790 100
rect 755 50 790 80
rect 755 30 765 50
rect 785 30 790 50
rect 755 20 790 30
rect 830 190 865 200
rect 830 170 835 190
rect 855 170 865 190
rect 830 140 865 170
rect 830 120 835 140
rect 855 120 865 140
rect 830 100 865 120
rect 830 80 835 100
rect 855 80 865 100
rect 830 50 865 80
rect 830 30 835 50
rect 855 30 865 50
rect 830 20 865 30
rect 880 190 915 200
rect 880 170 890 190
rect 910 170 915 190
rect 880 140 915 170
rect 880 120 890 140
rect 910 120 915 140
rect 880 100 915 120
rect 880 80 890 100
rect 910 80 915 100
rect 880 50 915 80
rect 880 30 890 50
rect 910 30 915 50
rect 880 20 915 30
rect 955 190 990 200
rect 955 170 960 190
rect 980 170 990 190
rect 955 140 990 170
rect 955 120 960 140
rect 980 120 990 140
rect 955 100 990 120
rect 955 80 960 100
rect 980 80 990 100
rect 955 50 990 80
rect 955 30 960 50
rect 980 30 990 50
rect 955 20 990 30
rect 1005 190 1040 200
rect 1005 170 1015 190
rect 1035 170 1040 190
rect 1005 140 1040 170
rect 1005 120 1015 140
rect 1035 120 1040 140
rect 1005 100 1040 120
rect 1005 80 1015 100
rect 1035 80 1040 100
rect 1005 50 1040 80
rect 1005 30 1015 50
rect 1035 30 1040 50
rect 1005 20 1040 30
rect 1080 190 1115 220
rect 1080 170 1085 190
rect 1105 170 1115 190
rect 1080 140 1115 170
rect 1080 120 1085 140
rect 1105 120 1115 140
rect 1080 100 1115 120
rect 1080 80 1085 100
rect 1105 80 1115 100
rect 1080 50 1115 80
rect 1080 30 1085 50
rect 1105 30 1115 50
rect 1080 20 1115 30
rect 1130 280 1165 290
rect 1130 260 1140 280
rect 1160 260 1165 280
rect 1130 240 1165 260
rect 1130 220 1140 240
rect 1160 220 1165 240
rect 1130 190 1165 220
rect 1130 170 1140 190
rect 1160 170 1165 190
rect 1130 140 1165 170
rect 1130 120 1140 140
rect 1160 120 1165 140
rect 1130 100 1165 120
rect 1130 80 1140 100
rect 1160 80 1165 100
rect 1130 50 1165 80
rect 1130 30 1140 50
rect 1160 30 1165 50
rect 1130 20 1165 30
rect 1205 280 1240 290
rect 1205 260 1210 280
rect 1230 260 1240 280
rect 1205 240 1240 260
rect 1205 220 1210 240
rect 1230 220 1240 240
rect 1205 190 1240 220
rect 1205 170 1210 190
rect 1230 170 1240 190
rect 1205 140 1240 170
rect 1205 120 1210 140
rect 1230 120 1240 140
rect 1205 100 1240 120
rect 1205 80 1210 100
rect 1230 80 1240 100
rect 1205 50 1240 80
rect 1205 30 1210 50
rect 1230 30 1240 50
rect 1205 20 1240 30
rect 1255 280 1290 290
rect 1255 260 1265 280
rect 1285 260 1290 280
rect 1255 240 1290 260
rect 1255 220 1265 240
rect 1285 220 1290 240
rect 1255 190 1290 220
rect 1255 170 1265 190
rect 1285 170 1290 190
rect 1255 140 1290 170
rect 1255 120 1265 140
rect 1285 120 1290 140
rect 1255 100 1290 120
rect 1255 80 1265 100
rect 1285 80 1290 100
rect 1255 50 1290 80
rect 1255 30 1265 50
rect 1285 30 1290 50
rect 1255 20 1290 30
rect 1330 280 1365 290
rect 1330 260 1335 280
rect 1355 260 1365 280
rect 1330 240 1365 260
rect 1330 220 1335 240
rect 1355 220 1365 240
rect 1330 190 1365 220
rect 1330 170 1335 190
rect 1355 170 1365 190
rect 1330 140 1365 170
rect 1330 120 1335 140
rect 1355 120 1365 140
rect 1330 100 1365 120
rect 1330 80 1335 100
rect 1355 80 1365 100
rect 1330 50 1365 80
rect 1330 30 1335 50
rect 1355 30 1365 50
rect 1330 20 1365 30
rect 1380 280 1415 290
rect 1380 260 1390 280
rect 1410 260 1415 280
rect 1380 240 1415 260
rect 1380 220 1390 240
rect 1410 220 1415 240
rect 1380 190 1415 220
rect 1380 170 1390 190
rect 1410 170 1415 190
rect 1380 140 1415 170
rect 1380 120 1390 140
rect 1410 120 1415 140
rect 1380 100 1415 120
rect 1380 80 1390 100
rect 1410 80 1415 100
rect 1380 50 1415 80
rect 1380 30 1390 50
rect 1410 30 1415 50
rect 1380 20 1415 30
rect 1455 100 1490 110
rect 1455 80 1460 100
rect 1480 80 1490 100
rect 1455 50 1490 80
rect 1455 30 1460 50
rect 1480 30 1490 50
rect 1455 20 1490 30
rect 1505 100 1540 110
rect 1505 80 1515 100
rect 1535 80 1540 100
rect 1505 50 1540 80
rect 1505 30 1515 50
rect 1535 30 1540 50
rect 1505 20 1540 30
rect 1595 100 1630 110
rect 1595 80 1600 100
rect 1620 80 1630 100
rect 1595 50 1630 80
rect 1595 30 1600 50
rect 1620 30 1630 50
rect 1595 20 1630 30
rect 1645 100 1680 110
rect 1645 80 1655 100
rect 1675 80 1680 100
rect 1645 50 1680 80
rect 1645 30 1655 50
rect 1675 30 1680 50
rect 1645 20 1680 30
rect 1725 100 1760 110
rect 1725 80 1730 100
rect 1750 80 1760 100
rect 1725 50 1760 80
rect 1725 30 1730 50
rect 1750 30 1760 50
rect 1725 20 1760 30
rect 1775 100 1810 110
rect 1775 80 1785 100
rect 1805 80 1810 100
rect 1775 50 1810 80
rect 1775 30 1785 50
rect 1805 30 1810 50
rect 1775 20 1810 30
rect 1850 100 1885 110
rect 1850 80 1855 100
rect 1875 80 1885 100
rect 1850 50 1885 80
rect 1850 30 1855 50
rect 1875 30 1885 50
rect 1850 20 1885 30
rect 1900 100 1935 110
rect 1900 80 1910 100
rect 1930 80 1935 100
rect 1900 50 1935 80
rect 1900 30 1910 50
rect 1930 30 1935 50
rect 1900 20 1935 30
<< ndiffc >>
rect -40 -205 -20 -185
rect -40 -255 -20 -235
rect 15 -205 35 -185
rect 15 -255 35 -235
rect 85 -205 105 -185
rect 85 -255 105 -235
rect 140 -205 160 -185
rect 140 -255 160 -235
rect 210 -205 230 -185
rect 210 -255 230 -235
rect 265 -205 285 -185
rect 265 -255 285 -235
rect 335 -205 355 -185
rect 335 -255 355 -235
rect 390 -205 410 -185
rect 390 -255 410 -235
rect 460 -205 480 -185
rect 460 -255 480 -235
rect 515 -205 535 -185
rect 515 -255 535 -235
rect 585 -205 605 -185
rect 585 -255 605 -235
rect 640 -205 660 -185
rect 640 -255 660 -235
rect 710 -205 730 -185
rect 710 -255 730 -235
rect 765 -205 785 -185
rect 765 -255 785 -235
rect 835 -205 855 -185
rect 835 -255 855 -235
rect 890 -205 910 -185
rect 890 -255 910 -235
rect 960 -205 980 -185
rect 960 -255 980 -235
rect 1015 -205 1035 -185
rect 1015 -255 1035 -235
rect 1085 -205 1105 -185
rect 1085 -255 1105 -235
rect 1085 -300 1105 -280
rect 1140 -205 1160 -185
rect 1140 -255 1160 -235
rect 1140 -300 1160 -280
rect 1210 -205 1230 -185
rect 1210 -255 1230 -235
rect 1210 -300 1230 -280
rect 1265 -205 1285 -185
rect 1265 -255 1285 -235
rect 1265 -300 1285 -280
rect 1335 -205 1355 -185
rect 1335 -255 1355 -235
rect 1335 -300 1355 -280
rect 1390 -205 1410 -185
rect 1460 -210 1480 -185
rect 1515 -210 1535 -185
rect 1600 -210 1620 -185
rect 1655 -210 1675 -185
rect 1730 -210 1750 -185
rect 1785 -210 1805 -185
rect 1855 -210 1875 -185
rect 1910 -210 1930 -185
rect 1390 -255 1410 -235
rect 1390 -300 1410 -280
<< pdiffc >>
rect 1085 260 1105 280
rect 1085 220 1105 240
rect -40 170 -20 190
rect -40 120 -20 140
rect -40 80 -20 100
rect -40 30 -20 50
rect 15 170 35 190
rect 15 120 35 140
rect 15 80 35 100
rect 15 30 35 50
rect 85 170 105 190
rect 85 120 105 140
rect 85 80 105 100
rect 85 30 105 50
rect 140 170 160 190
rect 140 120 160 140
rect 140 80 160 100
rect 140 30 160 50
rect 210 170 230 190
rect 210 120 230 140
rect 210 80 230 100
rect 210 30 230 50
rect 265 170 285 190
rect 265 120 285 140
rect 265 80 285 100
rect 265 30 285 50
rect 335 170 355 190
rect 335 120 355 140
rect 335 80 355 100
rect 335 30 355 50
rect 390 170 410 190
rect 390 120 410 140
rect 390 80 410 100
rect 390 30 410 50
rect 460 170 480 190
rect 460 120 480 140
rect 460 80 480 100
rect 460 30 480 50
rect 515 170 535 190
rect 515 120 535 140
rect 515 80 535 100
rect 515 30 535 50
rect 585 170 605 190
rect 585 120 605 140
rect 585 80 605 100
rect 585 30 605 50
rect 640 170 660 190
rect 640 120 660 140
rect 640 80 660 100
rect 640 30 660 50
rect 710 170 730 190
rect 710 120 730 140
rect 710 80 730 100
rect 710 30 730 50
rect 765 170 785 190
rect 765 120 785 140
rect 765 80 785 100
rect 765 30 785 50
rect 835 170 855 190
rect 835 120 855 140
rect 835 80 855 100
rect 835 30 855 50
rect 890 170 910 190
rect 890 120 910 140
rect 890 80 910 100
rect 890 30 910 50
rect 960 170 980 190
rect 960 120 980 140
rect 960 80 980 100
rect 960 30 980 50
rect 1015 170 1035 190
rect 1015 120 1035 140
rect 1015 80 1035 100
rect 1015 30 1035 50
rect 1085 170 1105 190
rect 1085 120 1105 140
rect 1085 80 1105 100
rect 1085 30 1105 50
rect 1140 260 1160 280
rect 1140 220 1160 240
rect 1140 170 1160 190
rect 1140 120 1160 140
rect 1140 80 1160 100
rect 1140 30 1160 50
rect 1210 260 1230 280
rect 1210 220 1230 240
rect 1210 170 1230 190
rect 1210 120 1230 140
rect 1210 80 1230 100
rect 1210 30 1230 50
rect 1265 260 1285 280
rect 1265 220 1285 240
rect 1265 170 1285 190
rect 1265 120 1285 140
rect 1265 80 1285 100
rect 1265 30 1285 50
rect 1335 260 1355 280
rect 1335 220 1355 240
rect 1335 170 1355 190
rect 1335 120 1355 140
rect 1335 80 1355 100
rect 1335 30 1355 50
rect 1390 260 1410 280
rect 1390 220 1410 240
rect 1390 170 1410 190
rect 1390 120 1410 140
rect 1390 80 1410 100
rect 1390 30 1410 50
rect 1460 80 1480 100
rect 1460 30 1480 50
rect 1515 80 1535 100
rect 1515 30 1535 50
rect 1600 80 1620 100
rect 1600 30 1620 50
rect 1655 80 1675 100
rect 1655 30 1675 50
rect 1730 80 1750 100
rect 1730 30 1750 50
rect 1785 80 1805 100
rect 1785 30 1805 50
rect 1855 80 1875 100
rect 1855 30 1875 50
rect 1910 80 1930 100
rect 1910 30 1930 50
<< psubdiff >>
rect 1450 -285 1545 -280
rect 1450 -305 1465 -285
rect 1485 -305 1510 -285
rect 1530 -305 1545 -285
rect 1450 -310 1545 -305
rect 1590 -285 1685 -280
rect 1590 -305 1605 -285
rect 1625 -305 1650 -285
rect 1670 -305 1685 -285
rect 1590 -310 1685 -305
rect 1720 -285 1815 -280
rect 1720 -305 1735 -285
rect 1755 -305 1780 -285
rect 1800 -305 1815 -285
rect 1720 -310 1815 -305
rect 1845 -285 1940 -280
rect 1845 -305 1860 -285
rect 1880 -305 1905 -285
rect 1925 -305 1940 -285
rect 1845 -310 1940 -305
rect -50 -330 45 -325
rect -50 -350 -35 -330
rect -15 -350 10 -330
rect 30 -350 45 -330
rect -50 -355 45 -350
rect 75 -330 170 -325
rect 75 -350 90 -330
rect 110 -350 135 -330
rect 155 -350 170 -330
rect 75 -355 170 -350
rect 200 -330 295 -325
rect 200 -350 215 -330
rect 235 -350 260 -330
rect 280 -350 295 -330
rect 200 -355 295 -350
rect 325 -330 420 -325
rect 325 -350 340 -330
rect 360 -350 385 -330
rect 405 -350 420 -330
rect 325 -355 420 -350
rect 450 -330 545 -325
rect 450 -350 465 -330
rect 485 -350 510 -330
rect 530 -350 545 -330
rect 450 -355 545 -350
rect 575 -330 670 -325
rect 575 -350 590 -330
rect 610 -350 635 -330
rect 655 -350 670 -330
rect 575 -355 670 -350
rect 700 -330 795 -325
rect 700 -350 715 -330
rect 735 -350 760 -330
rect 780 -350 795 -330
rect 700 -355 795 -350
rect 825 -330 920 -325
rect 825 -350 840 -330
rect 860 -350 885 -330
rect 905 -350 920 -330
rect 825 -355 920 -350
rect 950 -330 1045 -325
rect 950 -350 965 -330
rect 985 -350 1010 -330
rect 1030 -350 1045 -330
rect 950 -355 1045 -350
rect 1075 -360 1170 -355
rect 1075 -380 1090 -360
rect 1110 -380 1135 -360
rect 1155 -380 1170 -360
rect 1075 -385 1170 -380
rect 1200 -360 1295 -355
rect 1200 -380 1215 -360
rect 1235 -380 1260 -360
rect 1280 -380 1295 -360
rect 1200 -385 1295 -380
rect 1325 -360 1420 -355
rect 1325 -380 1340 -360
rect 1360 -380 1385 -360
rect 1405 -380 1420 -360
rect 1325 -385 1420 -380
<< nsubdiff >>
rect 1075 435 1170 440
rect 1075 415 1090 435
rect 1110 415 1135 435
rect 1155 415 1170 435
rect 1075 410 1170 415
rect 1200 435 1295 440
rect 1200 415 1215 435
rect 1235 415 1260 435
rect 1280 415 1295 435
rect 1200 410 1295 415
rect 1325 435 1420 440
rect 1325 415 1340 435
rect 1360 415 1385 435
rect 1405 415 1420 435
rect 1325 410 1420 415
rect -50 265 45 270
rect -50 245 -35 265
rect -15 245 10 265
rect 30 245 45 265
rect -50 240 45 245
rect 75 265 170 270
rect 75 245 90 265
rect 110 245 135 265
rect 155 245 170 265
rect 75 240 170 245
rect 200 265 295 270
rect 200 245 215 265
rect 235 245 260 265
rect 280 245 295 265
rect 200 240 295 245
rect 325 265 420 270
rect 325 245 340 265
rect 360 245 385 265
rect 405 245 420 265
rect 325 240 420 245
rect 450 265 545 270
rect 450 245 465 265
rect 485 245 510 265
rect 530 245 545 265
rect 450 240 545 245
rect 575 265 670 270
rect 575 245 590 265
rect 610 245 635 265
rect 655 245 670 265
rect 575 240 670 245
rect 700 265 795 270
rect 700 245 715 265
rect 735 245 760 265
rect 780 245 795 265
rect 700 240 795 245
rect 825 265 920 270
rect 825 245 840 265
rect 860 245 885 265
rect 905 245 920 265
rect 825 240 920 245
rect 950 265 1045 270
rect 950 245 965 265
rect 985 245 1010 265
rect 1030 245 1045 265
rect 950 240 1045 245
rect -40 230 -20 240
rect 585 230 605 240
rect 1450 170 1545 175
rect 1450 150 1465 170
rect 1485 150 1510 170
rect 1530 150 1545 170
rect 1450 145 1545 150
rect 1590 170 1685 175
rect 1590 150 1605 170
rect 1625 150 1650 170
rect 1670 150 1685 170
rect 1590 145 1685 150
rect 1720 170 1815 175
rect 1720 150 1735 170
rect 1755 150 1780 170
rect 1800 150 1815 170
rect 1720 145 1815 150
rect 1845 170 1940 175
rect 1845 150 1860 170
rect 1880 150 1905 170
rect 1925 150 1940 170
rect 1845 145 1940 150
<< psubdiffcont >>
rect 1465 -305 1485 -285
rect 1510 -305 1530 -285
rect 1605 -305 1625 -285
rect 1650 -305 1670 -285
rect 1735 -305 1755 -285
rect 1780 -305 1800 -285
rect 1860 -305 1880 -285
rect 1905 -305 1925 -285
rect -35 -350 -15 -330
rect 10 -350 30 -330
rect 90 -350 110 -330
rect 135 -350 155 -330
rect 215 -350 235 -330
rect 260 -350 280 -330
rect 340 -350 360 -330
rect 385 -350 405 -330
rect 465 -350 485 -330
rect 510 -350 530 -330
rect 590 -350 610 -330
rect 635 -350 655 -330
rect 715 -350 735 -330
rect 760 -350 780 -330
rect 840 -350 860 -330
rect 885 -350 905 -330
rect 965 -350 985 -330
rect 1010 -350 1030 -330
rect 1090 -380 1110 -360
rect 1135 -380 1155 -360
rect 1215 -380 1235 -360
rect 1260 -380 1280 -360
rect 1340 -380 1360 -360
rect 1385 -380 1405 -360
<< nsubdiffcont >>
rect 1090 415 1110 435
rect 1135 415 1155 435
rect 1215 415 1235 435
rect 1260 415 1280 435
rect 1340 415 1360 435
rect 1385 415 1405 435
rect -35 245 -15 265
rect 10 245 30 265
rect 90 245 110 265
rect 135 245 155 265
rect 215 245 235 265
rect 260 245 280 265
rect 340 245 360 265
rect 385 245 405 265
rect 465 245 485 265
rect 510 245 530 265
rect 590 245 610 265
rect 635 245 655 265
rect 715 245 735 265
rect 760 245 780 265
rect 840 245 860 265
rect 885 245 905 265
rect 965 245 985 265
rect 1010 245 1030 265
rect 1465 150 1485 170
rect 1510 150 1530 170
rect 1605 150 1625 170
rect 1650 150 1670 170
rect 1735 150 1755 170
rect 1780 150 1800 170
rect 1860 150 1880 170
rect 1905 150 1925 170
<< poly >>
rect 1115 290 1130 305
rect 1240 290 1255 305
rect 1365 290 1380 305
rect -10 200 5 215
rect 115 200 130 215
rect 240 200 255 215
rect 365 200 380 215
rect 490 200 505 215
rect 615 200 630 215
rect 740 200 755 215
rect 865 200 880 215
rect 990 200 1005 215
rect 1490 110 1505 125
rect 1630 110 1645 125
rect 1760 110 1775 125
rect 1885 110 1900 125
rect -10 -40 5 20
rect 115 -40 130 20
rect 240 -40 255 20
rect 365 -40 380 20
rect 490 -40 505 20
rect 615 -40 630 20
rect 740 -40 755 20
rect 865 -40 880 20
rect 990 -40 1005 20
rect -10 -45 30 -40
rect -10 -65 0 -45
rect 20 -65 30 -45
rect -10 -70 30 -65
rect 115 -45 155 -40
rect 115 -65 125 -45
rect 145 -65 155 -45
rect 115 -70 155 -65
rect 240 -45 280 -40
rect 240 -65 250 -45
rect 270 -65 280 -45
rect 240 -70 280 -65
rect 365 -45 405 -40
rect 365 -65 375 -45
rect 395 -65 405 -45
rect 365 -70 405 -65
rect 490 -45 530 -40
rect 490 -65 500 -45
rect 520 -65 530 -45
rect 490 -70 530 -65
rect 615 -45 655 -40
rect 615 -65 625 -45
rect 645 -65 655 -45
rect 615 -70 655 -65
rect 740 -45 780 -40
rect 740 -65 750 -45
rect 770 -65 780 -45
rect 740 -70 780 -65
rect 865 -45 905 -40
rect 865 -65 875 -45
rect 895 -65 905 -45
rect 865 -70 905 -65
rect 965 -45 1005 -40
rect 965 -65 975 -45
rect 995 -65 1005 -45
rect 965 -70 1005 -65
rect -10 -175 5 -70
rect 115 -175 130 -70
rect 240 -175 255 -70
rect 365 -175 380 -70
rect 490 -175 505 -70
rect 615 -175 630 -70
rect 740 -175 755 -70
rect 865 -175 880 -70
rect 990 -175 1005 -70
rect 1115 -40 1130 20
rect 1240 -40 1255 20
rect 1365 -40 1380 20
rect 1115 -45 1155 -40
rect 1115 -65 1125 -45
rect 1145 -65 1155 -45
rect 1115 -70 1155 -65
rect 1240 -45 1280 -40
rect 1240 -65 1250 -45
rect 1270 -65 1280 -45
rect 1240 -70 1280 -65
rect 1335 -45 1380 -40
rect 1335 -65 1345 -45
rect 1365 -65 1380 -45
rect 1335 -70 1380 -65
rect 1115 -175 1130 -70
rect 1240 -175 1255 -70
rect 1365 -175 1380 -70
rect 1490 -90 1505 20
rect 1630 -90 1645 20
rect 1760 -15 1775 20
rect 1725 -20 1775 -15
rect 1725 -40 1735 -20
rect 1755 -40 1775 -20
rect 1725 -45 1775 -40
rect 1465 -95 1505 -90
rect 1465 -115 1475 -95
rect 1495 -115 1505 -95
rect 1465 -120 1505 -115
rect 1605 -95 1645 -90
rect 1605 -115 1615 -95
rect 1635 -115 1645 -95
rect 1605 -120 1645 -115
rect 1490 -175 1505 -120
rect 1630 -175 1645 -120
rect 1760 -175 1775 -45
rect 1885 -50 1900 20
rect 1850 -55 1900 -50
rect 1850 -75 1860 -55
rect 1880 -75 1900 -55
rect 1850 -80 1900 -75
rect 1885 -175 1900 -80
rect -10 -280 5 -265
rect 115 -280 130 -265
rect 240 -280 255 -265
rect 365 -280 380 -265
rect 490 -280 505 -265
rect 615 -280 630 -265
rect 740 -280 755 -265
rect 865 -280 880 -265
rect 990 -280 1005 -265
rect 1490 -235 1505 -220
rect 1630 -235 1645 -220
rect 1760 -235 1775 -220
rect 1885 -235 1900 -220
rect 1115 -325 1130 -310
rect 1240 -325 1255 -310
rect 1365 -325 1380 -310
<< polycont >>
rect 0 -65 20 -45
rect 125 -65 145 -45
rect 250 -65 270 -45
rect 375 -65 395 -45
rect 500 -65 520 -45
rect 625 -65 645 -45
rect 750 -65 770 -45
rect 875 -65 895 -45
rect 975 -65 995 -45
rect 1125 -65 1145 -45
rect 1250 -65 1270 -45
rect 1345 -65 1365 -45
rect 1735 -40 1755 -20
rect 1475 -115 1495 -95
rect 1615 -115 1635 -95
rect 1860 -75 1880 -55
<< locali >>
rect 1075 435 1170 440
rect 1075 415 1090 435
rect 1110 415 1130 435
rect 1155 415 1170 435
rect 1075 410 1170 415
rect 1200 435 1295 440
rect 1200 415 1215 435
rect 1235 415 1255 435
rect 1280 415 1295 435
rect 1200 410 1295 415
rect 1325 435 1420 440
rect 1325 415 1340 435
rect 1360 415 1380 435
rect 1405 415 1420 435
rect 1325 410 1420 415
rect 1085 290 1105 410
rect 1080 280 1110 290
rect -50 265 45 270
rect -50 245 -35 265
rect -15 245 5 265
rect 30 245 45 265
rect -50 240 45 245
rect 75 265 170 270
rect 75 245 90 265
rect 110 245 130 265
rect 155 245 170 265
rect 75 240 170 245
rect 200 265 295 270
rect 200 245 215 265
rect 235 245 255 265
rect 280 245 295 265
rect 200 240 295 245
rect 325 265 420 270
rect 325 245 340 265
rect 360 245 380 265
rect 405 245 420 265
rect 325 240 420 245
rect 450 265 545 270
rect 450 245 465 265
rect 485 245 505 265
rect 530 245 545 265
rect 450 240 545 245
rect 575 265 670 270
rect 575 245 590 265
rect 610 245 630 265
rect 655 245 670 265
rect 575 240 670 245
rect 700 265 795 270
rect 700 245 715 265
rect 735 245 755 265
rect 780 245 795 265
rect 700 240 795 245
rect 825 265 920 270
rect 825 245 840 265
rect 860 245 880 265
rect 905 245 920 265
rect 825 240 920 245
rect 950 265 1045 270
rect 950 245 965 265
rect 985 245 1005 265
rect 1030 245 1045 265
rect 950 240 1045 245
rect 1080 260 1085 280
rect 1105 260 1110 280
rect 1080 240 1110 260
rect -40 200 -20 240
rect 85 200 105 240
rect 335 200 355 240
rect 585 200 605 240
rect 710 200 730 240
rect 835 200 855 240
rect 1080 220 1085 240
rect 1105 220 1110 240
rect -45 190 -15 200
rect -45 170 -40 190
rect -20 170 -15 190
rect -45 140 -15 170
rect -45 120 -40 140
rect -20 120 -15 140
rect -45 100 -15 120
rect -45 80 -40 100
rect -20 80 -15 100
rect -45 50 -15 80
rect -45 30 -40 50
rect -20 30 -15 50
rect -45 20 -15 30
rect 10 190 40 200
rect 10 170 15 190
rect 35 170 40 190
rect 10 140 40 170
rect 10 120 15 140
rect 35 120 40 140
rect 10 100 40 120
rect 10 80 15 100
rect 35 80 40 100
rect 10 50 40 80
rect 10 30 15 50
rect 35 30 40 50
rect 10 20 40 30
rect 80 190 110 200
rect 80 170 85 190
rect 105 170 110 190
rect 80 140 110 170
rect 80 120 85 140
rect 105 120 110 140
rect 80 100 110 120
rect 80 80 85 100
rect 105 80 110 100
rect 80 50 110 80
rect 80 30 85 50
rect 105 30 110 50
rect 80 20 110 30
rect 135 190 165 200
rect 135 170 140 190
rect 160 170 165 190
rect 135 140 165 170
rect 135 120 140 140
rect 160 120 165 140
rect 135 100 165 120
rect 135 80 140 100
rect 160 80 165 100
rect 135 50 165 80
rect 135 30 140 50
rect 160 30 165 50
rect 135 20 165 30
rect 205 190 235 200
rect 205 170 210 190
rect 230 170 235 190
rect 205 140 235 170
rect 205 120 210 140
rect 230 120 235 140
rect 205 100 235 120
rect 205 80 210 100
rect 230 80 235 100
rect 205 50 235 80
rect 205 30 210 50
rect 230 30 235 50
rect 205 20 235 30
rect 260 190 290 200
rect 260 170 265 190
rect 285 170 290 190
rect 260 140 290 170
rect 260 120 265 140
rect 285 120 290 140
rect 260 100 290 120
rect 260 80 265 100
rect 285 80 290 100
rect 260 50 290 80
rect 260 30 265 50
rect 285 30 290 50
rect 260 20 290 30
rect 330 190 360 200
rect 330 170 335 190
rect 355 170 360 190
rect 330 140 360 170
rect 330 120 335 140
rect 355 120 360 140
rect 330 100 360 120
rect 330 80 335 100
rect 355 80 360 100
rect 330 50 360 80
rect 330 30 335 50
rect 355 30 360 50
rect 330 20 360 30
rect 385 190 415 200
rect 385 170 390 190
rect 410 170 415 190
rect 385 140 415 170
rect 385 120 390 140
rect 410 120 415 140
rect 385 100 415 120
rect 385 80 390 100
rect 410 80 415 100
rect 385 50 415 80
rect 385 30 390 50
rect 410 30 415 50
rect 385 20 415 30
rect 455 190 485 200
rect 455 170 460 190
rect 480 170 485 190
rect 455 140 485 170
rect 455 120 460 140
rect 480 120 485 140
rect 455 100 485 120
rect 455 80 460 100
rect 480 80 485 100
rect 455 50 485 80
rect 455 30 460 50
rect 480 30 485 50
rect 455 20 485 30
rect 510 190 540 200
rect 510 170 515 190
rect 535 170 540 190
rect 510 140 540 170
rect 510 120 515 140
rect 535 120 540 140
rect 510 100 540 120
rect 510 80 515 100
rect 535 80 540 100
rect 510 50 540 80
rect 510 30 515 50
rect 535 30 540 50
rect 510 20 540 30
rect 580 190 610 200
rect 580 170 585 190
rect 605 170 610 190
rect 580 140 610 170
rect 580 120 585 140
rect 605 120 610 140
rect 580 100 610 120
rect 580 80 585 100
rect 605 80 610 100
rect 580 50 610 80
rect 580 30 585 50
rect 605 30 610 50
rect 580 20 610 30
rect 635 190 665 200
rect 635 170 640 190
rect 660 170 665 190
rect 635 140 665 170
rect 635 120 640 140
rect 660 120 665 140
rect 635 100 665 120
rect 635 80 640 100
rect 660 80 665 100
rect 635 50 665 80
rect 635 30 640 50
rect 660 30 665 50
rect 635 20 665 30
rect 705 190 735 200
rect 705 170 710 190
rect 730 170 735 190
rect 705 140 735 170
rect 705 120 710 140
rect 730 120 735 140
rect 705 100 735 120
rect 705 80 710 100
rect 730 80 735 100
rect 705 50 735 80
rect 705 30 710 50
rect 730 30 735 50
rect 705 20 735 30
rect 760 190 790 200
rect 760 170 765 190
rect 785 170 790 190
rect 760 140 790 170
rect 760 120 765 140
rect 785 120 790 140
rect 760 100 790 120
rect 760 80 765 100
rect 785 80 790 100
rect 760 50 790 80
rect 760 30 765 50
rect 785 30 790 50
rect 760 20 790 30
rect 830 190 860 200
rect 830 170 835 190
rect 855 170 860 190
rect 830 140 860 170
rect 830 120 835 140
rect 855 120 860 140
rect 830 100 860 120
rect 830 80 835 100
rect 855 80 860 100
rect 830 50 860 80
rect 830 30 835 50
rect 855 30 860 50
rect 830 20 860 30
rect 885 190 915 200
rect 885 170 890 190
rect 910 170 915 190
rect 885 140 915 170
rect 885 120 890 140
rect 910 120 915 140
rect 885 100 915 120
rect 885 80 890 100
rect 910 80 915 100
rect 885 50 915 80
rect 885 30 890 50
rect 910 30 915 50
rect 885 20 915 30
rect 955 190 985 200
rect 955 170 960 190
rect 980 170 985 190
rect 955 140 985 170
rect 955 120 960 140
rect 980 120 985 140
rect 955 100 985 120
rect 955 80 960 100
rect 980 80 985 100
rect 955 50 985 80
rect 955 30 960 50
rect 980 30 985 50
rect 955 20 985 30
rect 1010 190 1040 200
rect 1010 170 1015 190
rect 1035 170 1040 190
rect 1010 140 1040 170
rect 1010 120 1015 140
rect 1035 120 1040 140
rect 1010 100 1040 120
rect 1010 80 1015 100
rect 1035 80 1040 100
rect 1010 50 1040 80
rect 1010 30 1015 50
rect 1035 30 1040 50
rect 1010 20 1040 30
rect 1080 190 1110 220
rect 1080 170 1085 190
rect 1105 170 1110 190
rect 1080 140 1110 170
rect 1080 120 1085 140
rect 1105 120 1110 140
rect 1080 100 1110 120
rect 1080 80 1085 100
rect 1105 80 1110 100
rect 1080 50 1110 80
rect 1080 30 1085 50
rect 1105 30 1110 50
rect 1080 20 1110 30
rect 1135 280 1165 290
rect 1135 260 1140 280
rect 1160 260 1165 280
rect 1135 240 1165 260
rect 1135 220 1140 240
rect 1160 220 1165 240
rect 1135 190 1165 220
rect 1135 170 1140 190
rect 1160 170 1165 190
rect 1135 140 1165 170
rect 1135 120 1140 140
rect 1160 120 1165 140
rect 1135 100 1165 120
rect 1135 80 1140 100
rect 1160 80 1165 100
rect 1135 50 1165 80
rect 1135 30 1140 50
rect 1160 30 1165 50
rect 1135 20 1165 30
rect 1205 280 1235 290
rect 1205 260 1210 280
rect 1230 260 1235 280
rect 1205 240 1235 260
rect 1205 220 1210 240
rect 1230 220 1235 240
rect 1205 190 1235 220
rect 1205 170 1210 190
rect 1230 170 1235 190
rect 1205 140 1235 170
rect 1205 120 1210 140
rect 1230 120 1235 140
rect 1205 100 1235 120
rect 1205 80 1210 100
rect 1230 80 1235 100
rect 1205 50 1235 80
rect 1205 30 1210 50
rect 1230 30 1235 50
rect 1205 20 1235 30
rect 1260 280 1290 290
rect 1260 260 1265 280
rect 1285 260 1290 280
rect 1260 240 1290 260
rect 1260 220 1265 240
rect 1285 220 1290 240
rect 1260 190 1290 220
rect 1260 170 1265 190
rect 1285 170 1290 190
rect 1260 140 1290 170
rect 1260 120 1265 140
rect 1285 120 1290 140
rect 1260 100 1290 120
rect 1260 80 1265 100
rect 1285 80 1290 100
rect 1260 50 1290 80
rect 1260 30 1265 50
rect 1285 30 1290 50
rect 1260 20 1290 30
rect 1330 280 1360 290
rect 1330 260 1335 280
rect 1355 260 1360 280
rect 1330 240 1360 260
rect 1330 220 1335 240
rect 1355 220 1360 240
rect 1330 190 1360 220
rect 1330 170 1335 190
rect 1355 170 1360 190
rect 1330 140 1360 170
rect 1330 120 1335 140
rect 1355 120 1360 140
rect 1330 100 1360 120
rect 1330 80 1335 100
rect 1355 80 1360 100
rect 1330 50 1360 80
rect 1330 30 1335 50
rect 1355 30 1360 50
rect 1330 20 1360 30
rect 1385 280 1415 290
rect 1385 260 1390 280
rect 1410 260 1415 280
rect 1385 240 1415 260
rect 1385 220 1390 240
rect 1410 220 1415 240
rect 1385 190 1415 220
rect 1385 170 1390 190
rect 1410 170 1415 190
rect 1385 140 1415 170
rect 1450 170 1545 175
rect 1450 150 1465 170
rect 1485 150 1510 170
rect 1530 150 1545 170
rect 1450 145 1545 150
rect 1590 170 1685 175
rect 1590 150 1605 170
rect 1625 150 1650 170
rect 1670 150 1685 170
rect 1590 145 1685 150
rect 1720 170 1815 175
rect 1720 150 1735 170
rect 1755 150 1780 170
rect 1800 150 1815 170
rect 1720 145 1815 150
rect 1845 170 1940 175
rect 1845 150 1860 170
rect 1880 150 1905 170
rect 1925 150 1940 170
rect 1845 145 1940 150
rect 1385 120 1390 140
rect 1410 120 1415 140
rect 1385 100 1415 120
rect 1460 110 1480 145
rect 1600 110 1620 145
rect 1730 110 1750 145
rect 1855 110 1875 145
rect 1385 80 1390 100
rect 1410 80 1415 100
rect 1385 50 1415 80
rect 1385 30 1390 50
rect 1410 30 1415 50
rect 1385 20 1415 30
rect 1455 100 1485 110
rect 1455 80 1460 100
rect 1480 80 1485 100
rect 1455 50 1485 80
rect 1455 30 1460 50
rect 1480 30 1485 50
rect 1455 20 1485 30
rect 1510 100 1560 110
rect 1510 80 1515 100
rect 1535 80 1560 100
rect 1510 50 1560 80
rect 1510 30 1515 50
rect 1535 30 1560 50
rect 1510 20 1560 30
rect 1595 100 1625 110
rect 1595 80 1600 100
rect 1620 80 1625 100
rect 1595 50 1625 80
rect 1595 30 1600 50
rect 1620 30 1625 50
rect 1595 20 1625 30
rect 1650 100 1700 110
rect 1650 80 1655 100
rect 1675 80 1700 100
rect 1650 50 1700 80
rect 1650 30 1655 50
rect 1675 30 1700 50
rect 1650 20 1700 30
rect 1725 100 1755 110
rect 1725 80 1730 100
rect 1750 80 1755 100
rect 1725 50 1755 80
rect 1725 30 1730 50
rect 1750 30 1755 50
rect 1725 20 1755 30
rect 1780 100 1810 110
rect 1780 80 1785 100
rect 1805 80 1810 100
rect 1780 50 1810 80
rect 1780 30 1785 50
rect 1805 30 1810 50
rect 1780 20 1810 30
rect 1850 100 1880 110
rect 1850 80 1855 100
rect 1875 80 1880 100
rect 1850 50 1880 80
rect 1850 30 1855 50
rect 1875 30 1880 50
rect 1850 20 1880 30
rect 1905 100 1935 110
rect 1905 80 1910 100
rect 1930 80 1935 100
rect 1905 50 1935 80
rect 1905 30 1910 50
rect 1930 30 1935 50
rect 1905 20 1935 30
rect 15 0 35 20
rect 140 0 160 20
rect 210 0 230 20
rect 15 -20 230 0
rect 265 0 285 20
rect 390 0 410 20
rect 460 0 480 20
rect 265 -20 320 0
rect 390 -20 480 0
rect 515 0 535 20
rect 640 0 660 20
rect 765 0 785 20
rect 890 0 910 20
rect 960 0 980 20
rect 515 -20 570 0
rect 640 -20 980 0
rect 1015 0 1035 20
rect 1140 0 1160 20
rect 1210 0 1230 20
rect 1015 -20 1070 0
rect 1140 -20 1230 0
rect 1265 0 1285 20
rect 1335 0 1355 20
rect 1265 -20 1355 0
rect 1390 0 1410 20
rect 1390 -20 1420 0
rect -10 -45 30 -40
rect -10 -65 0 -45
rect 20 -65 30 -45
rect -10 -70 30 -65
rect 115 -45 155 -40
rect 115 -65 125 -45
rect 145 -65 155 -45
rect 115 -70 155 -65
rect 240 -45 280 -40
rect 240 -65 250 -45
rect 270 -65 280 -45
rect 240 -70 280 -65
rect 300 -95 320 -20
rect 365 -45 405 -40
rect 365 -65 375 -45
rect 395 -65 405 -45
rect 365 -70 405 -65
rect 490 -45 530 -40
rect 490 -65 500 -45
rect 520 -65 530 -45
rect 490 -70 530 -65
rect 550 -85 570 -20
rect 615 -45 655 -40
rect 615 -65 625 -45
rect 645 -65 655 -45
rect 615 -70 655 -65
rect 740 -45 780 -40
rect 740 -65 750 -45
rect 770 -65 780 -45
rect 740 -70 780 -65
rect 865 -45 905 -40
rect 865 -65 875 -45
rect 895 -65 905 -45
rect 865 -70 905 -65
rect 965 -45 1005 -40
rect 965 -65 975 -45
rect 995 -65 1005 -45
rect 965 -70 1005 -65
rect 540 -90 580 -85
rect 540 -95 550 -90
rect 15 -115 230 -95
rect 15 -175 35 -115
rect 140 -175 160 -115
rect 210 -175 230 -115
rect 265 -110 550 -95
rect 570 -95 580 -90
rect 965 -95 985 -70
rect 1050 -95 1070 -20
rect 1115 -45 1155 -40
rect 1115 -65 1125 -45
rect 1145 -65 1155 -45
rect 1115 -70 1155 -65
rect 1240 -45 1280 -40
rect 1240 -65 1250 -45
rect 1270 -65 1280 -45
rect 1240 -70 1280 -65
rect 1335 -45 1375 -40
rect 1335 -65 1345 -45
rect 1365 -65 1375 -45
rect 1335 -70 1375 -65
rect 1400 -95 1420 -20
rect 1540 -15 1560 20
rect 1540 -20 1580 -15
rect 1540 -40 1550 -20
rect 1570 -40 1580 -20
rect 1540 -45 1580 -40
rect 1465 -95 1505 -90
rect 570 -110 985 -95
rect 265 -115 985 -110
rect 1015 -115 1475 -95
rect 1495 -115 1505 -95
rect 265 -175 285 -115
rect 515 -175 535 -115
rect 640 -155 980 -135
rect 640 -175 660 -155
rect 765 -175 785 -155
rect 890 -175 910 -155
rect 960 -175 980 -155
rect 1015 -175 1035 -115
rect 1140 -155 1230 -135
rect 1140 -175 1160 -155
rect 1210 -175 1230 -155
rect 1265 -155 1355 -135
rect 1265 -175 1285 -155
rect 1335 -175 1355 -155
rect 1390 -175 1410 -115
rect 1465 -120 1505 -115
rect 1540 -175 1560 -45
rect 1680 -90 1700 20
rect 1725 -20 1765 -15
rect 1725 -40 1735 -20
rect 1755 -40 1765 -20
rect 1725 -45 1765 -40
rect 1790 -55 1810 20
rect 1910 -50 1930 20
rect 1850 -55 1890 -50
rect 1790 -75 1860 -55
rect 1880 -75 1890 -55
rect 1605 -95 1645 -90
rect 1605 -115 1615 -95
rect 1635 -115 1645 -95
rect 1605 -120 1645 -115
rect 1680 -95 1720 -90
rect 1680 -115 1690 -95
rect 1710 -115 1720 -95
rect 1680 -120 1720 -115
rect 1680 -175 1700 -120
rect 1790 -175 1810 -75
rect 1850 -80 1890 -75
rect 1910 -55 1960 -50
rect 1910 -75 1930 -55
rect 1950 -75 1960 -55
rect 1910 -80 1960 -75
rect 1910 -175 1930 -80
rect -45 -185 -15 -175
rect -45 -205 -40 -185
rect -20 -205 -15 -185
rect -45 -235 -15 -205
rect -45 -255 -40 -235
rect -20 -255 -15 -235
rect -45 -265 -15 -255
rect 10 -185 40 -175
rect 10 -205 15 -185
rect 35 -205 40 -185
rect 10 -235 40 -205
rect 10 -255 15 -235
rect 35 -255 40 -235
rect 10 -265 40 -255
rect 80 -185 110 -175
rect 80 -205 85 -185
rect 105 -205 110 -185
rect 80 -235 110 -205
rect 80 -255 85 -235
rect 105 -255 110 -235
rect 80 -265 110 -255
rect 135 -185 165 -175
rect 135 -205 140 -185
rect 160 -205 165 -185
rect 135 -235 165 -205
rect 135 -255 140 -235
rect 160 -255 165 -235
rect 135 -265 165 -255
rect 205 -185 235 -175
rect 205 -205 210 -185
rect 230 -205 235 -185
rect 205 -235 235 -205
rect 205 -255 210 -235
rect 230 -255 235 -235
rect 205 -265 235 -255
rect 260 -185 290 -175
rect 260 -205 265 -185
rect 285 -205 290 -185
rect 260 -235 290 -205
rect 260 -255 265 -235
rect 285 -255 290 -235
rect 260 -265 290 -255
rect 330 -185 360 -175
rect 330 -205 335 -185
rect 355 -205 360 -185
rect 330 -235 360 -205
rect 330 -255 335 -235
rect 355 -255 360 -235
rect 330 -265 360 -255
rect 385 -185 415 -175
rect 385 -205 390 -185
rect 410 -205 415 -185
rect 385 -235 415 -205
rect 385 -255 390 -235
rect 410 -255 415 -235
rect 385 -265 415 -255
rect 455 -185 485 -175
rect 455 -205 460 -185
rect 480 -205 485 -185
rect 455 -235 485 -205
rect 455 -255 460 -235
rect 480 -255 485 -235
rect 455 -265 485 -255
rect 510 -185 540 -175
rect 510 -205 515 -185
rect 535 -205 540 -185
rect 510 -235 540 -205
rect 510 -255 515 -235
rect 535 -255 540 -235
rect 510 -265 540 -255
rect 580 -185 610 -175
rect 580 -205 585 -185
rect 605 -205 610 -185
rect 580 -235 610 -205
rect 580 -255 585 -235
rect 605 -255 610 -235
rect 580 -265 610 -255
rect 635 -185 665 -175
rect 635 -205 640 -185
rect 660 -205 665 -185
rect 635 -235 665 -205
rect 635 -255 640 -235
rect 660 -255 665 -235
rect 635 -265 665 -255
rect 705 -185 735 -175
rect 705 -205 710 -185
rect 730 -205 735 -185
rect 705 -235 735 -205
rect 705 -255 710 -235
rect 730 -255 735 -235
rect 705 -265 735 -255
rect 760 -185 790 -175
rect 760 -205 765 -185
rect 785 -205 790 -185
rect 760 -235 790 -205
rect 760 -255 765 -235
rect 785 -255 790 -235
rect 760 -265 790 -255
rect 830 -185 860 -175
rect 830 -205 835 -185
rect 855 -205 860 -185
rect 830 -235 860 -205
rect 830 -255 835 -235
rect 855 -255 860 -235
rect 830 -265 860 -255
rect 885 -185 915 -175
rect 885 -205 890 -185
rect 910 -205 915 -185
rect 885 -235 915 -205
rect 885 -255 890 -235
rect 910 -255 915 -235
rect 885 -265 915 -255
rect 955 -185 985 -175
rect 955 -205 960 -185
rect 980 -205 985 -185
rect 955 -235 985 -205
rect 955 -255 960 -235
rect 980 -255 985 -235
rect 955 -265 985 -255
rect 1010 -185 1040 -175
rect 1010 -205 1015 -185
rect 1035 -205 1040 -185
rect 1010 -235 1040 -205
rect 1010 -255 1015 -235
rect 1035 -255 1040 -235
rect 1010 -265 1040 -255
rect 1080 -185 1110 -175
rect 1080 -205 1085 -185
rect 1105 -205 1110 -185
rect 1080 -235 1110 -205
rect 1080 -255 1085 -235
rect 1105 -255 1110 -235
rect -40 -325 -20 -265
rect 85 -325 105 -265
rect 335 -325 355 -265
rect 390 -285 410 -265
rect 460 -285 480 -265
rect 390 -305 480 -285
rect 585 -325 605 -265
rect 710 -325 730 -265
rect 835 -325 855 -265
rect 1080 -280 1110 -255
rect 1080 -300 1085 -280
rect 1105 -300 1110 -280
rect 1080 -310 1110 -300
rect 1135 -185 1165 -175
rect 1135 -205 1140 -185
rect 1160 -205 1165 -185
rect 1135 -235 1165 -205
rect 1135 -255 1140 -235
rect 1160 -255 1165 -235
rect 1135 -280 1165 -255
rect 1135 -300 1140 -280
rect 1160 -300 1165 -280
rect 1135 -310 1165 -300
rect 1205 -185 1235 -175
rect 1205 -205 1210 -185
rect 1230 -205 1235 -185
rect 1205 -235 1235 -205
rect 1205 -255 1210 -235
rect 1230 -255 1235 -235
rect 1205 -280 1235 -255
rect 1205 -300 1210 -280
rect 1230 -300 1235 -280
rect 1205 -310 1235 -300
rect 1260 -185 1290 -175
rect 1260 -205 1265 -185
rect 1285 -205 1290 -185
rect 1260 -235 1290 -205
rect 1260 -255 1265 -235
rect 1285 -255 1290 -235
rect 1260 -280 1290 -255
rect 1260 -300 1265 -280
rect 1285 -300 1290 -280
rect 1260 -310 1290 -300
rect 1330 -185 1360 -175
rect 1330 -205 1335 -185
rect 1355 -205 1360 -185
rect 1330 -235 1360 -205
rect 1330 -255 1335 -235
rect 1355 -255 1360 -235
rect 1330 -280 1360 -255
rect 1330 -300 1335 -280
rect 1355 -300 1360 -280
rect 1330 -310 1360 -300
rect 1385 -185 1415 -175
rect 1385 -205 1390 -185
rect 1410 -205 1415 -185
rect 1385 -235 1415 -205
rect 1455 -185 1485 -175
rect 1455 -210 1460 -185
rect 1480 -210 1485 -185
rect 1455 -220 1485 -210
rect 1510 -185 1560 -175
rect 1510 -210 1515 -185
rect 1535 -210 1560 -185
rect 1510 -220 1560 -210
rect 1595 -185 1625 -175
rect 1595 -210 1600 -185
rect 1620 -210 1625 -185
rect 1595 -220 1625 -210
rect 1650 -185 1700 -175
rect 1650 -210 1655 -185
rect 1675 -210 1700 -185
rect 1650 -220 1700 -210
rect 1725 -185 1755 -175
rect 1725 -210 1730 -185
rect 1750 -210 1755 -185
rect 1725 -220 1755 -210
rect 1780 -185 1810 -175
rect 1780 -210 1785 -185
rect 1805 -210 1810 -185
rect 1780 -220 1810 -210
rect 1850 -185 1880 -175
rect 1850 -210 1855 -185
rect 1875 -210 1880 -185
rect 1850 -220 1880 -210
rect 1905 -185 1935 -175
rect 1905 -210 1910 -185
rect 1930 -210 1935 -185
rect 1905 -220 1935 -210
rect 1385 -255 1390 -235
rect 1410 -255 1415 -235
rect 1385 -280 1415 -255
rect 1460 -280 1480 -220
rect 1600 -280 1620 -220
rect 1730 -280 1750 -220
rect 1855 -280 1875 -220
rect 1385 -300 1390 -280
rect 1410 -300 1415 -280
rect 1385 -310 1415 -300
rect 1450 -285 1545 -280
rect 1450 -305 1465 -285
rect 1485 -305 1510 -285
rect 1530 -305 1545 -285
rect 1450 -310 1545 -305
rect 1590 -285 1685 -280
rect 1590 -305 1605 -285
rect 1625 -305 1650 -285
rect 1670 -305 1685 -285
rect 1590 -310 1685 -305
rect 1720 -285 1815 -280
rect 1720 -305 1735 -285
rect 1755 -305 1780 -285
rect 1800 -305 1815 -285
rect 1720 -310 1815 -305
rect 1845 -285 1940 -280
rect 1845 -305 1860 -285
rect 1880 -305 1905 -285
rect 1925 -305 1940 -285
rect 1845 -310 1940 -305
rect -50 -330 45 -325
rect -50 -350 -35 -330
rect -15 -350 10 -330
rect 30 -350 45 -330
rect -50 -355 45 -350
rect 75 -330 170 -325
rect 75 -350 90 -330
rect 110 -350 135 -330
rect 155 -350 170 -330
rect 75 -355 170 -350
rect 200 -330 295 -325
rect 200 -350 215 -330
rect 235 -350 260 -330
rect 280 -350 295 -330
rect 200 -355 295 -350
rect 325 -330 420 -325
rect 325 -350 340 -330
rect 360 -350 385 -330
rect 405 -350 420 -330
rect 325 -355 420 -350
rect 450 -330 545 -325
rect 450 -350 465 -330
rect 485 -350 510 -330
rect 530 -350 545 -330
rect 450 -355 545 -350
rect 575 -330 670 -325
rect 575 -350 590 -330
rect 610 -350 635 -330
rect 655 -350 670 -330
rect 575 -355 670 -350
rect 700 -330 795 -325
rect 700 -350 715 -330
rect 735 -350 760 -330
rect 780 -350 795 -330
rect 700 -355 795 -350
rect 825 -330 920 -325
rect 825 -350 840 -330
rect 860 -350 885 -330
rect 905 -350 920 -330
rect 825 -355 920 -350
rect 950 -330 1045 -325
rect 950 -350 965 -330
rect 985 -350 1010 -330
rect 1030 -350 1045 -330
rect 950 -355 1045 -350
rect 1085 -355 1105 -310
rect 1075 -360 1170 -355
rect 1075 -380 1090 -360
rect 1110 -380 1135 -360
rect 1155 -380 1170 -360
rect 1075 -385 1170 -380
rect 1200 -360 1295 -355
rect 1200 -380 1215 -360
rect 1235 -380 1260 -360
rect 1280 -380 1295 -360
rect 1200 -385 1295 -380
rect 1325 -360 1420 -355
rect 1325 -380 1340 -360
rect 1360 -380 1385 -360
rect 1405 -380 1420 -360
rect 1325 -385 1420 -380
<< viali >>
rect 1130 415 1135 435
rect 1135 415 1150 435
rect 1255 415 1260 435
rect 1260 415 1275 435
rect 1380 415 1385 435
rect 1385 415 1400 435
rect 5 245 10 265
rect 10 245 25 265
rect 130 245 135 265
rect 135 245 150 265
rect 255 245 260 265
rect 260 245 275 265
rect 380 245 385 265
rect 385 245 400 265
rect 505 245 510 265
rect 510 245 525 265
rect 630 245 635 265
rect 635 245 650 265
rect 755 245 760 265
rect 760 245 775 265
rect 880 245 885 265
rect 885 245 900 265
rect 1005 245 1010 265
rect 1010 245 1025 265
rect 1510 150 1530 170
rect 1650 150 1670 170
rect 1780 150 1800 170
rect 1905 150 1925 170
rect 0 -65 20 -45
rect 125 -65 145 -45
rect 250 -65 270 -45
rect 375 -65 395 -45
rect 500 -65 520 -45
rect 625 -65 645 -45
rect 750 -65 770 -45
rect 875 -65 895 -45
rect 550 -110 570 -90
rect 1125 -65 1145 -45
rect 1250 -65 1270 -45
rect 1345 -65 1365 -45
rect 1550 -40 1570 -20
rect 1735 -40 1755 -20
rect 1615 -115 1635 -95
rect 1690 -115 1710 -95
rect 1930 -75 1950 -55
rect 1510 -305 1530 -285
rect 1650 -305 1670 -285
rect 1780 -305 1800 -285
rect 1905 -305 1925 -285
rect 10 -350 30 -330
rect 135 -350 155 -330
rect 260 -350 280 -330
rect 385 -350 405 -330
rect 510 -350 530 -330
rect 635 -350 655 -330
rect 760 -350 780 -330
rect 885 -350 905 -330
rect 1010 -350 1030 -330
rect 1135 -380 1155 -360
rect 1260 -380 1280 -360
rect 1385 -380 1405 -360
<< metal1 >>
rect -85 475 1925 495
rect 5 270 25 475
rect 40 340 80 345
rect 40 310 45 340
rect 75 310 80 340
rect 40 305 80 310
rect -5 265 35 270
rect -5 245 5 265
rect 25 245 35 265
rect -5 240 35 245
rect 50 -40 70 305
rect 130 270 150 475
rect 165 390 205 395
rect 165 360 170 390
rect 200 360 205 390
rect 165 355 205 360
rect 120 265 160 270
rect 120 245 130 265
rect 150 245 160 265
rect 120 240 160 245
rect 175 -40 195 355
rect 255 270 275 475
rect 290 440 330 445
rect 290 410 295 440
rect 325 410 330 440
rect 290 405 330 410
rect 245 265 285 270
rect 245 245 255 265
rect 275 245 285 265
rect 245 240 285 245
rect 300 -40 320 405
rect 380 270 400 475
rect 415 390 455 395
rect 415 360 420 390
rect 450 360 455 390
rect 415 355 455 360
rect 370 265 410 270
rect 370 245 380 265
rect 400 245 410 265
rect 370 240 410 245
rect 425 -40 445 355
rect 505 270 525 475
rect 540 340 580 345
rect 540 310 545 340
rect 575 310 580 340
rect 540 305 580 310
rect 495 265 535 270
rect 495 245 505 265
rect 525 245 535 265
rect 495 240 535 245
rect 550 -40 570 305
rect 630 270 650 475
rect 665 340 705 345
rect 665 310 670 340
rect 700 310 705 340
rect 665 305 705 310
rect 620 265 660 270
rect 620 245 630 265
rect 650 245 660 265
rect 620 240 660 245
rect 675 -40 695 305
rect 755 270 775 475
rect 790 390 830 395
rect 790 360 795 390
rect 825 360 830 390
rect 790 355 830 360
rect 745 265 785 270
rect 745 245 755 265
rect 775 245 785 265
rect 745 240 785 245
rect 800 -40 820 355
rect 880 270 900 475
rect 915 440 955 445
rect 915 410 920 440
rect 950 410 955 440
rect 915 405 955 410
rect 870 265 910 270
rect 870 245 880 265
rect 900 245 910 265
rect 870 240 910 245
rect 925 -40 945 405
rect 1005 270 1025 475
rect 1130 440 1150 475
rect 1255 440 1275 475
rect 1380 440 1400 475
rect 1445 440 1485 445
rect 1120 435 1160 440
rect 1120 415 1130 435
rect 1150 415 1160 435
rect 1120 410 1160 415
rect 1245 435 1285 440
rect 1245 415 1255 435
rect 1275 415 1285 435
rect 1245 410 1285 415
rect 1370 435 1410 440
rect 1370 415 1380 435
rect 1400 415 1410 435
rect 1370 410 1410 415
rect 1445 410 1450 440
rect 1480 410 1485 440
rect 1445 405 1485 410
rect 1290 390 1330 395
rect 1290 360 1295 390
rect 1325 360 1330 390
rect 1455 375 1475 405
rect 1290 355 1330 360
rect 1425 355 1475 375
rect 1165 340 1205 345
rect 1165 310 1170 340
rect 1200 310 1205 340
rect 1165 305 1205 310
rect 995 265 1035 270
rect 995 245 1005 265
rect 1025 245 1035 265
rect 995 240 1035 245
rect 1175 -40 1195 305
rect 1300 -40 1320 355
rect -10 -45 70 -40
rect -10 -65 0 -45
rect 20 -65 70 -45
rect -10 -70 70 -65
rect 115 -45 195 -40
rect 115 -65 125 -45
rect 145 -65 195 -45
rect 115 -70 195 -65
rect 240 -45 320 -40
rect 240 -65 250 -45
rect 270 -65 320 -45
rect 240 -70 320 -65
rect 365 -45 445 -40
rect 365 -65 375 -45
rect 395 -65 445 -45
rect 365 -70 445 -65
rect 490 -45 570 -40
rect 490 -65 500 -45
rect 520 -65 570 -45
rect 490 -70 570 -65
rect 615 -45 695 -40
rect 615 -65 625 -45
rect 645 -65 695 -45
rect 615 -70 695 -65
rect 740 -45 820 -40
rect 740 -65 750 -45
rect 770 -65 820 -45
rect 740 -70 820 -65
rect 865 -45 945 -40
rect 865 -65 875 -45
rect 895 -65 945 -45
rect 865 -70 945 -65
rect 1115 -45 1195 -40
rect 1115 -65 1125 -45
rect 1145 -65 1195 -45
rect 1115 -70 1195 -65
rect 1240 -45 1320 -40
rect 1240 -65 1250 -45
rect 1270 -65 1320 -45
rect 1240 -70 1320 -65
rect 1335 -45 1375 -40
rect 1425 -45 1445 355
rect 1510 175 1530 475
rect 1650 175 1670 475
rect 1780 175 1800 475
rect 1905 175 1925 475
rect 1500 170 1540 175
rect 1500 150 1510 170
rect 1530 150 1540 170
rect 1500 145 1540 150
rect 1640 170 1680 175
rect 1640 150 1650 170
rect 1670 150 1680 170
rect 1640 145 1680 150
rect 1770 170 1810 175
rect 1770 150 1780 170
rect 1800 150 1810 170
rect 1770 145 1810 150
rect 1895 170 1935 175
rect 1895 150 1905 170
rect 1925 150 1935 170
rect 1895 145 1935 150
rect 1540 -20 1580 -15
rect 1725 -20 1765 -15
rect 1540 -40 1550 -20
rect 1570 -40 1735 -20
rect 1755 -40 1765 -20
rect 1540 -45 1580 -40
rect 1725 -45 1765 -40
rect 1335 -65 1345 -45
rect 1365 -65 1445 -45
rect 1920 -55 1960 -50
rect 1335 -70 1375 -65
rect 1920 -75 1930 -55
rect 1950 -75 2000 -55
rect 1920 -80 1960 -75
rect 540 -90 580 -85
rect 540 -110 550 -90
rect 570 -110 580 -90
rect 1605 -95 1645 -90
rect 540 -115 580 -110
rect 1585 -115 1615 -95
rect 1635 -115 1645 -95
rect 550 -295 570 -115
rect 1585 -120 1645 -115
rect 1680 -95 1720 -90
rect 1680 -115 1690 -95
rect 1710 -115 2000 -95
rect 1680 -120 1720 -115
rect 1585 -140 1605 -120
rect 1425 -160 1605 -140
rect 1425 -295 1445 -160
rect 550 -310 1445 -295
rect 1500 -285 1540 -280
rect 1500 -305 1510 -285
rect 1530 -305 1540 -285
rect 1500 -310 1540 -305
rect 1640 -285 1680 -280
rect 1640 -305 1650 -285
rect 1670 -305 1680 -285
rect 1640 -310 1680 -305
rect 1770 -285 1810 -280
rect 1770 -305 1780 -285
rect 1800 -305 1810 -285
rect 1770 -310 1810 -305
rect 1895 -285 1935 -280
rect 1895 -305 1905 -285
rect 1925 -305 1935 -285
rect 1895 -310 1935 -305
rect 0 -330 40 -325
rect 0 -350 10 -330
rect 30 -350 40 -330
rect 0 -355 40 -350
rect 125 -330 165 -325
rect 125 -350 135 -330
rect 155 -350 165 -330
rect 125 -355 165 -350
rect 250 -330 290 -325
rect 250 -350 260 -330
rect 280 -350 290 -330
rect 250 -355 290 -350
rect 375 -330 415 -325
rect 375 -350 385 -330
rect 405 -350 415 -330
rect 375 -355 415 -350
rect 500 -330 540 -325
rect 500 -350 510 -330
rect 530 -350 540 -330
rect 500 -355 540 -350
rect 625 -330 665 -325
rect 625 -350 635 -330
rect 655 -350 665 -330
rect 625 -355 665 -350
rect 750 -330 790 -325
rect 750 -350 760 -330
rect 780 -350 790 -330
rect 750 -355 790 -350
rect 875 -330 915 -325
rect 875 -350 885 -330
rect 905 -350 915 -330
rect 875 -355 915 -350
rect 1000 -330 1040 -325
rect 1000 -350 1010 -330
rect 1030 -350 1040 -330
rect 1000 -355 1040 -350
rect 10 -440 30 -355
rect 135 -440 155 -355
rect 260 -440 280 -355
rect 385 -440 405 -355
rect 510 -440 530 -355
rect 635 -440 655 -355
rect 760 -440 780 -355
rect 885 -440 905 -355
rect 1010 -440 1030 -355
rect 1125 -360 1165 -355
rect 1125 -380 1135 -360
rect 1155 -380 1165 -360
rect 1125 -385 1165 -380
rect 1250 -360 1290 -355
rect 1250 -380 1260 -360
rect 1280 -380 1290 -360
rect 1250 -385 1290 -380
rect 1375 -360 1415 -355
rect 1375 -380 1385 -360
rect 1405 -380 1415 -360
rect 1375 -385 1415 -380
rect 1135 -440 1155 -385
rect 1260 -440 1280 -385
rect 1385 -440 1405 -385
rect 1510 -440 1530 -310
rect 1650 -440 1670 -310
rect 1780 -440 1800 -310
rect 1905 -440 1925 -310
rect -90 -460 1925 -440
<< via1 >>
rect 45 310 75 340
rect 170 360 200 390
rect 295 410 325 440
rect 420 360 450 390
rect 545 310 575 340
rect 670 310 700 340
rect 795 360 825 390
rect 920 410 950 440
rect 1450 410 1480 440
rect 1295 360 1325 390
rect 1170 310 1200 340
<< metal2 >>
rect 290 440 330 445
rect 290 435 295 440
rect -85 415 295 435
rect 290 410 295 415
rect 325 435 330 440
rect 915 440 955 445
rect 915 435 920 440
rect 325 415 920 435
rect 325 410 330 415
rect 290 405 330 410
rect 915 410 920 415
rect 950 435 955 440
rect 1445 440 1485 445
rect 1445 435 1450 440
rect 950 415 1450 435
rect 950 410 955 415
rect 915 405 955 410
rect 1445 410 1450 415
rect 1480 410 1485 440
rect 1445 405 1485 410
rect 165 390 205 395
rect 165 385 170 390
rect -85 365 170 385
rect 165 360 170 365
rect 200 385 205 390
rect 415 390 455 395
rect 415 385 420 390
rect 200 365 420 385
rect 200 360 205 365
rect 165 355 205 360
rect 415 360 420 365
rect 450 385 455 390
rect 790 390 830 395
rect 790 385 795 390
rect 450 365 795 385
rect 450 360 455 365
rect 415 355 455 360
rect 790 360 795 365
rect 825 385 830 390
rect 1290 390 1330 395
rect 1290 385 1295 390
rect 825 365 1295 385
rect 825 360 830 365
rect 790 355 830 360
rect 1290 360 1295 365
rect 1325 360 1330 390
rect 1290 355 1330 360
rect 40 340 80 345
rect 40 335 45 340
rect -85 315 45 335
rect 40 310 45 315
rect 75 335 80 340
rect 540 340 580 345
rect 540 335 545 340
rect 75 315 545 335
rect 75 310 80 315
rect 40 305 80 310
rect 540 310 545 315
rect 575 335 580 340
rect 665 340 705 345
rect 665 335 670 340
rect 575 315 670 335
rect 575 310 580 315
rect 540 305 580 310
rect 665 310 670 315
rect 700 335 705 340
rect 1165 340 1205 345
rect 1165 335 1170 340
rect 700 315 1170 335
rect 700 310 705 315
rect 665 305 705 310
rect 1165 310 1170 315
rect 1200 310 1205 340
rect 1165 305 1205 310
<< labels >>
rlabel metal2 -65 315 -55 335 1 a
rlabel metal2 -65 365 -55 385 1 b
rlabel metal2 -65 415 -55 435 1 cin
rlabel metal1 -60 485 -60 485 1 vdd
rlabel metal1 -50 -455 -50 -455 1 gnd
rlabel metal1 1985 -75 1995 -55 1 sum
rlabel metal1 1985 -115 1995 -95 1 cout
<< end >>
