magic
tech sky130A
timestamp 1720937323
<< nwell >>
rect 1180 440 1990 690
rect 1335 410 1990 440
<< nmos >>
rect 1240 320 1255 365
rect 1915 300 1930 345
rect 1395 170 1410 260
rect 1520 170 1535 260
rect 1645 170 1660 260
rect 1770 170 1785 260
<< pmos >>
rect 1240 460 1255 550
rect 1395 430 1410 610
rect 1520 430 1535 610
rect 1645 430 1660 610
rect 1770 430 1785 610
rect 1915 440 1930 530
<< ndiff >>
rect 1205 355 1240 365
rect 1205 330 1210 355
rect 1230 330 1240 355
rect 1205 320 1240 330
rect 1255 355 1290 365
rect 1255 330 1265 355
rect 1285 330 1290 355
rect 1255 320 1290 330
rect 1880 335 1915 345
rect 1880 310 1885 335
rect 1905 310 1915 335
rect 1880 300 1915 310
rect 1930 335 1965 345
rect 1930 310 1940 335
rect 1960 310 1965 335
rect 1930 300 1965 310
rect 1360 250 1395 260
rect 1360 230 1365 250
rect 1385 230 1395 250
rect 1360 200 1395 230
rect 1360 180 1365 200
rect 1385 180 1395 200
rect 1360 170 1395 180
rect 1410 250 1445 260
rect 1410 230 1420 250
rect 1440 230 1445 250
rect 1410 200 1445 230
rect 1410 180 1420 200
rect 1440 180 1445 200
rect 1410 170 1445 180
rect 1485 250 1520 260
rect 1485 230 1490 250
rect 1510 230 1520 250
rect 1485 200 1520 230
rect 1485 180 1490 200
rect 1510 180 1520 200
rect 1485 170 1520 180
rect 1535 250 1570 260
rect 1535 230 1545 250
rect 1565 230 1570 250
rect 1535 200 1570 230
rect 1535 180 1545 200
rect 1565 180 1570 200
rect 1535 170 1570 180
rect 1610 250 1645 260
rect 1610 230 1615 250
rect 1635 230 1645 250
rect 1610 200 1645 230
rect 1610 180 1615 200
rect 1635 180 1645 200
rect 1610 170 1645 180
rect 1660 250 1695 260
rect 1660 230 1670 250
rect 1690 230 1695 250
rect 1660 200 1695 230
rect 1660 180 1670 200
rect 1690 180 1695 200
rect 1660 170 1695 180
rect 1735 250 1770 260
rect 1735 230 1740 250
rect 1760 230 1770 250
rect 1735 200 1770 230
rect 1735 180 1740 200
rect 1760 180 1770 200
rect 1735 170 1770 180
rect 1785 250 1820 260
rect 1785 230 1795 250
rect 1815 230 1820 250
rect 1785 200 1820 230
rect 1785 180 1795 200
rect 1815 180 1820 200
rect 1785 170 1820 180
<< pdiff >>
rect 1360 600 1395 610
rect 1360 580 1365 600
rect 1385 580 1395 600
rect 1360 560 1395 580
rect 1205 540 1240 550
rect 1205 520 1210 540
rect 1230 520 1240 540
rect 1205 490 1240 520
rect 1205 470 1210 490
rect 1230 470 1240 490
rect 1205 460 1240 470
rect 1255 540 1290 550
rect 1255 520 1265 540
rect 1285 520 1290 540
rect 1255 490 1290 520
rect 1255 470 1265 490
rect 1285 470 1290 490
rect 1255 460 1290 470
rect 1360 540 1365 560
rect 1385 540 1395 560
rect 1360 500 1395 540
rect 1360 480 1365 500
rect 1385 480 1395 500
rect 1360 460 1395 480
rect 1360 440 1365 460
rect 1385 440 1395 460
rect 1360 430 1395 440
rect 1410 600 1445 610
rect 1410 580 1420 600
rect 1440 580 1445 600
rect 1410 560 1445 580
rect 1410 540 1420 560
rect 1440 540 1445 560
rect 1410 500 1445 540
rect 1410 480 1420 500
rect 1440 480 1445 500
rect 1410 460 1445 480
rect 1410 440 1420 460
rect 1440 440 1445 460
rect 1410 430 1445 440
rect 1485 600 1520 610
rect 1485 580 1490 600
rect 1510 580 1520 600
rect 1485 560 1520 580
rect 1485 540 1490 560
rect 1510 540 1520 560
rect 1485 500 1520 540
rect 1485 480 1490 500
rect 1510 480 1520 500
rect 1485 460 1520 480
rect 1485 440 1490 460
rect 1510 440 1520 460
rect 1485 430 1520 440
rect 1535 600 1570 610
rect 1535 580 1545 600
rect 1565 580 1570 600
rect 1535 560 1570 580
rect 1535 540 1545 560
rect 1565 540 1570 560
rect 1535 500 1570 540
rect 1535 480 1545 500
rect 1565 480 1570 500
rect 1535 460 1570 480
rect 1535 440 1545 460
rect 1565 440 1570 460
rect 1535 430 1570 440
rect 1610 600 1645 610
rect 1610 580 1615 600
rect 1635 580 1645 600
rect 1610 560 1645 580
rect 1610 540 1615 560
rect 1635 540 1645 560
rect 1610 500 1645 540
rect 1610 480 1615 500
rect 1635 480 1645 500
rect 1610 460 1645 480
rect 1610 440 1615 460
rect 1635 440 1645 460
rect 1610 430 1645 440
rect 1660 600 1695 610
rect 1660 580 1670 600
rect 1690 580 1695 600
rect 1660 560 1695 580
rect 1660 540 1670 560
rect 1690 540 1695 560
rect 1660 500 1695 540
rect 1660 480 1670 500
rect 1690 480 1695 500
rect 1660 460 1695 480
rect 1660 440 1670 460
rect 1690 440 1695 460
rect 1660 430 1695 440
rect 1735 600 1770 610
rect 1735 580 1740 600
rect 1760 580 1770 600
rect 1735 560 1770 580
rect 1735 540 1740 560
rect 1760 540 1770 560
rect 1735 500 1770 540
rect 1735 480 1740 500
rect 1760 480 1770 500
rect 1735 460 1770 480
rect 1735 440 1740 460
rect 1760 440 1770 460
rect 1735 430 1770 440
rect 1785 600 1820 610
rect 1785 580 1795 600
rect 1815 580 1820 600
rect 1785 560 1820 580
rect 1785 540 1795 560
rect 1815 540 1820 560
rect 1785 500 1820 540
rect 1785 480 1795 500
rect 1815 480 1820 500
rect 1785 460 1820 480
rect 1785 440 1795 460
rect 1815 440 1820 460
rect 1880 520 1915 530
rect 1880 500 1885 520
rect 1905 500 1915 520
rect 1880 470 1915 500
rect 1880 450 1885 470
rect 1905 450 1915 470
rect 1880 440 1915 450
rect 1930 520 1965 530
rect 1930 500 1940 520
rect 1960 500 1965 520
rect 1930 470 1965 500
rect 1930 450 1940 470
rect 1960 450 1965 470
rect 1930 440 1965 450
rect 1785 430 1820 440
<< ndiffc >>
rect 1210 330 1230 355
rect 1265 330 1285 355
rect 1885 310 1905 335
rect 1940 310 1960 335
rect 1365 230 1385 250
rect 1365 180 1385 200
rect 1420 230 1440 250
rect 1420 180 1440 200
rect 1490 230 1510 250
rect 1490 180 1510 200
rect 1545 230 1565 250
rect 1545 180 1565 200
rect 1615 230 1635 250
rect 1615 180 1635 200
rect 1670 230 1690 250
rect 1670 180 1690 200
rect 1740 230 1760 250
rect 1740 180 1760 200
rect 1795 230 1815 250
rect 1795 180 1815 200
<< pdiffc >>
rect 1365 580 1385 600
rect 1210 520 1230 540
rect 1210 470 1230 490
rect 1265 520 1285 540
rect 1265 470 1285 490
rect 1365 540 1385 560
rect 1365 480 1385 500
rect 1365 440 1385 460
rect 1420 580 1440 600
rect 1420 540 1440 560
rect 1420 480 1440 500
rect 1420 440 1440 460
rect 1490 580 1510 600
rect 1490 540 1510 560
rect 1490 480 1510 500
rect 1490 440 1510 460
rect 1545 580 1565 600
rect 1545 540 1565 560
rect 1545 480 1565 500
rect 1545 440 1565 460
rect 1615 580 1635 600
rect 1615 540 1635 560
rect 1615 480 1635 500
rect 1615 440 1635 460
rect 1670 580 1690 600
rect 1670 540 1690 560
rect 1670 480 1690 500
rect 1670 440 1690 460
rect 1740 580 1760 600
rect 1740 540 1760 560
rect 1740 480 1760 500
rect 1740 440 1760 460
rect 1795 580 1815 600
rect 1795 540 1815 560
rect 1795 480 1815 500
rect 1795 440 1815 460
rect 1885 500 1905 520
rect 1885 450 1905 470
rect 1940 500 1960 520
rect 1940 450 1960 470
<< psubdiff >>
rect 1200 225 1295 230
rect 1200 205 1215 225
rect 1235 205 1260 225
rect 1280 205 1295 225
rect 1200 200 1295 205
rect 1875 205 1970 210
rect 1875 185 1890 205
rect 1910 185 1935 205
rect 1955 185 1970 205
rect 1875 180 1970 185
rect 1355 85 1450 90
rect 1355 65 1370 85
rect 1390 65 1415 85
rect 1435 65 1450 85
rect 1355 60 1450 65
rect 1480 85 1575 90
rect 1480 65 1495 85
rect 1515 65 1540 85
rect 1560 65 1575 85
rect 1480 60 1575 65
rect 1605 85 1700 90
rect 1605 65 1620 85
rect 1640 65 1665 85
rect 1685 65 1700 85
rect 1605 60 1700 65
rect 1730 85 1825 90
rect 1730 65 1745 85
rect 1765 65 1790 85
rect 1810 65 1825 85
rect 1730 60 1825 65
<< nsubdiff >>
rect 1355 665 1450 670
rect 1355 645 1370 665
rect 1390 645 1415 665
rect 1435 645 1450 665
rect 1355 640 1450 645
rect 1480 665 1575 670
rect 1480 645 1495 665
rect 1515 645 1540 665
rect 1560 645 1575 665
rect 1480 640 1575 645
rect 1605 665 1700 670
rect 1605 645 1620 665
rect 1640 645 1665 665
rect 1685 645 1700 665
rect 1605 640 1700 645
rect 1730 665 1825 670
rect 1730 645 1745 665
rect 1765 645 1790 665
rect 1810 645 1825 665
rect 1730 640 1825 645
rect 1200 605 1295 610
rect 1200 585 1215 605
rect 1235 585 1260 605
rect 1280 585 1295 605
rect 1200 580 1295 585
rect 1875 585 1970 590
rect 1875 565 1890 585
rect 1910 565 1935 585
rect 1955 565 1970 585
rect 1875 560 1970 565
<< psubdiffcont >>
rect 1215 205 1235 225
rect 1260 205 1280 225
rect 1890 185 1910 205
rect 1935 185 1955 205
rect 1370 65 1390 85
rect 1415 65 1435 85
rect 1495 65 1515 85
rect 1540 65 1560 85
rect 1620 65 1640 85
rect 1665 65 1685 85
rect 1745 65 1765 85
rect 1790 65 1810 85
<< nsubdiffcont >>
rect 1370 645 1390 665
rect 1415 645 1435 665
rect 1495 645 1515 665
rect 1540 645 1560 665
rect 1620 645 1640 665
rect 1665 645 1685 665
rect 1745 645 1765 665
rect 1790 645 1810 665
rect 1215 585 1235 605
rect 1260 585 1280 605
rect 1890 565 1910 585
rect 1935 565 1955 585
<< poly >>
rect 1395 610 1410 625
rect 1520 610 1535 625
rect 1645 610 1660 625
rect 1770 610 1785 625
rect 1240 550 1255 565
rect 1240 420 1255 460
rect 1915 530 1930 545
rect 1205 415 1255 420
rect 1205 395 1215 415
rect 1235 395 1255 415
rect 1205 390 1255 395
rect 1240 365 1255 390
rect 1395 360 1410 430
rect 1370 355 1410 360
rect 1520 355 1535 430
rect 1370 335 1380 355
rect 1400 335 1410 355
rect 1370 330 1410 335
rect 1240 305 1255 320
rect 1395 260 1410 330
rect 1495 350 1535 355
rect 1495 330 1505 350
rect 1525 330 1535 350
rect 1495 325 1535 330
rect 1520 260 1535 325
rect 1645 315 1660 430
rect 1620 310 1660 315
rect 1620 290 1630 310
rect 1650 290 1660 310
rect 1620 285 1660 290
rect 1645 260 1660 285
rect 1770 325 1785 430
rect 1915 400 1930 440
rect 1880 395 1930 400
rect 1880 375 1890 395
rect 1910 375 1930 395
rect 1880 370 1930 375
rect 1915 345 1930 370
rect 1770 315 1815 325
rect 1770 295 1785 315
rect 1805 295 1815 315
rect 1770 285 1815 295
rect 1915 285 1930 300
rect 1770 260 1785 285
rect 1395 155 1410 170
rect 1520 155 1535 170
rect 1645 155 1660 170
rect 1770 155 1785 170
<< polycont >>
rect 1215 395 1235 415
rect 1380 335 1400 355
rect 1505 330 1525 350
rect 1630 290 1650 310
rect 1890 375 1910 395
rect 1785 295 1805 315
<< locali >>
rect 1355 665 1450 670
rect 1355 645 1370 665
rect 1390 645 1415 665
rect 1435 645 1450 665
rect 1355 640 1450 645
rect 1480 665 1575 670
rect 1480 645 1495 665
rect 1515 645 1540 665
rect 1560 645 1575 665
rect 1480 640 1575 645
rect 1605 665 1700 670
rect 1605 645 1620 665
rect 1640 645 1665 665
rect 1685 645 1700 665
rect 1605 640 1700 645
rect 1730 665 1825 670
rect 1730 645 1745 665
rect 1765 645 1790 665
rect 1810 645 1825 665
rect 1730 640 1825 645
rect 1365 610 1385 640
rect 1490 610 1510 640
rect 1200 605 1295 610
rect 1200 585 1215 605
rect 1235 585 1260 605
rect 1280 585 1295 605
rect 1200 580 1295 585
rect 1360 600 1390 610
rect 1360 580 1365 600
rect 1385 580 1390 600
rect 1210 550 1230 580
rect 1360 560 1390 580
rect 1205 540 1235 550
rect 1205 520 1210 540
rect 1230 520 1235 540
rect 1205 490 1235 520
rect 1205 470 1210 490
rect 1230 470 1235 490
rect 1205 460 1235 470
rect 1260 540 1290 550
rect 1260 520 1265 540
rect 1285 520 1290 540
rect 1260 490 1290 520
rect 1260 470 1265 490
rect 1285 470 1290 490
rect 1260 460 1290 470
rect 1360 540 1365 560
rect 1385 540 1390 560
rect 1360 500 1390 540
rect 1360 480 1365 500
rect 1385 480 1390 500
rect 1360 460 1390 480
rect 1205 415 1245 420
rect 1205 395 1215 415
rect 1235 395 1245 415
rect 1205 390 1245 395
rect 1265 365 1285 460
rect 1360 440 1365 460
rect 1385 440 1390 460
rect 1360 430 1390 440
rect 1415 600 1445 610
rect 1415 580 1420 600
rect 1440 580 1445 600
rect 1415 560 1445 580
rect 1415 540 1420 560
rect 1440 540 1445 560
rect 1415 500 1445 540
rect 1415 480 1420 500
rect 1440 480 1445 500
rect 1415 460 1445 480
rect 1415 440 1420 460
rect 1440 440 1445 460
rect 1415 430 1445 440
rect 1485 600 1515 610
rect 1485 580 1490 600
rect 1510 580 1515 600
rect 1485 560 1515 580
rect 1485 540 1490 560
rect 1510 540 1515 560
rect 1485 500 1515 540
rect 1485 480 1490 500
rect 1510 480 1515 500
rect 1485 460 1515 480
rect 1485 440 1490 460
rect 1510 440 1515 460
rect 1485 430 1515 440
rect 1540 600 1570 610
rect 1540 580 1545 600
rect 1565 580 1570 600
rect 1540 560 1570 580
rect 1540 540 1545 560
rect 1565 540 1570 560
rect 1540 500 1570 540
rect 1540 480 1545 500
rect 1565 480 1570 500
rect 1540 460 1570 480
rect 1540 440 1545 460
rect 1565 440 1570 460
rect 1540 430 1570 440
rect 1610 600 1640 610
rect 1610 580 1615 600
rect 1635 580 1640 600
rect 1610 560 1640 580
rect 1610 540 1615 560
rect 1635 540 1640 560
rect 1610 500 1640 540
rect 1610 480 1615 500
rect 1635 480 1640 500
rect 1610 460 1640 480
rect 1610 440 1615 460
rect 1635 440 1640 460
rect 1610 430 1640 440
rect 1665 600 1695 610
rect 1665 580 1670 600
rect 1690 580 1695 600
rect 1665 560 1695 580
rect 1665 540 1670 560
rect 1690 540 1695 560
rect 1665 500 1695 540
rect 1665 480 1670 500
rect 1690 480 1695 500
rect 1665 460 1695 480
rect 1665 440 1670 460
rect 1690 440 1695 460
rect 1665 430 1695 440
rect 1735 600 1765 610
rect 1735 580 1740 600
rect 1760 580 1765 600
rect 1735 560 1765 580
rect 1735 540 1740 560
rect 1760 540 1765 560
rect 1735 500 1765 540
rect 1735 480 1740 500
rect 1760 480 1765 500
rect 1735 460 1765 480
rect 1735 440 1740 460
rect 1760 440 1765 460
rect 1735 430 1765 440
rect 1790 600 1820 610
rect 1790 580 1795 600
rect 1815 580 1820 600
rect 1790 560 1820 580
rect 1875 585 1970 590
rect 1875 565 1890 585
rect 1910 565 1935 585
rect 1955 565 1970 585
rect 1875 560 1970 565
rect 1790 540 1795 560
rect 1815 540 1820 560
rect 1790 500 1820 540
rect 1885 530 1905 560
rect 1790 480 1795 500
rect 1815 480 1820 500
rect 1790 460 1820 480
rect 1790 440 1795 460
rect 1815 440 1820 460
rect 1880 520 1910 530
rect 1880 500 1885 520
rect 1905 500 1910 520
rect 1880 470 1910 500
rect 1880 450 1885 470
rect 1905 450 1910 470
rect 1880 440 1910 450
rect 1935 520 1965 530
rect 1935 500 1940 520
rect 1960 500 1965 520
rect 1935 470 1965 500
rect 1935 450 1940 470
rect 1960 450 1965 470
rect 1935 440 1965 450
rect 1790 430 1820 440
rect 1420 405 1440 430
rect 1545 405 1565 430
rect 1615 405 1635 430
rect 1670 405 1690 430
rect 1420 385 1635 405
rect 1205 355 1235 365
rect 1205 330 1210 355
rect 1230 330 1235 355
rect 1205 320 1235 330
rect 1260 355 1290 365
rect 1260 330 1265 355
rect 1285 330 1290 355
rect 1370 355 1410 360
rect 1615 355 1635 385
rect 1660 400 1700 405
rect 1660 380 1670 400
rect 1690 380 1700 400
rect 1660 375 1700 380
rect 1740 355 1760 430
rect 1795 405 1815 430
rect 1785 400 1825 405
rect 1785 380 1795 400
rect 1815 380 1825 400
rect 1785 375 1825 380
rect 1880 395 1920 400
rect 1880 375 1890 395
rect 1910 375 1920 395
rect 1880 370 1920 375
rect 1370 335 1380 355
rect 1400 335 1410 355
rect 1370 330 1410 335
rect 1495 350 1535 355
rect 1495 330 1505 350
rect 1525 330 1535 350
rect 1615 335 1760 355
rect 1940 345 1960 440
rect 1880 335 1910 345
rect 1260 320 1290 330
rect 1495 325 1535 330
rect 1210 230 1230 320
rect 1265 300 1285 320
rect 1775 315 1815 325
rect 1620 310 1660 315
rect 1255 295 1295 300
rect 1255 275 1265 295
rect 1285 275 1295 295
rect 1620 290 1630 310
rect 1650 290 1660 310
rect 1620 285 1660 290
rect 1775 295 1785 315
rect 1805 295 1815 315
rect 1880 310 1885 335
rect 1905 310 1910 335
rect 1880 300 1910 310
rect 1935 335 1965 345
rect 1935 310 1940 335
rect 1960 310 1965 335
rect 1935 300 1965 310
rect 1775 285 1815 295
rect 1255 270 1295 275
rect 1360 250 1390 260
rect 1360 230 1365 250
rect 1385 230 1390 250
rect 1200 225 1295 230
rect 1200 205 1215 225
rect 1235 205 1260 225
rect 1280 205 1295 225
rect 1200 200 1295 205
rect 1360 200 1390 230
rect 1320 180 1365 200
rect 1385 180 1390 200
rect 1320 145 1340 180
rect 1360 170 1390 180
rect 1415 250 1445 260
rect 1415 230 1420 250
rect 1440 230 1445 250
rect 1415 200 1445 230
rect 1485 250 1515 260
rect 1485 230 1490 250
rect 1510 230 1515 250
rect 1485 200 1515 230
rect 1415 180 1420 200
rect 1440 180 1490 200
rect 1510 180 1515 200
rect 1415 170 1445 180
rect 1485 170 1515 180
rect 1540 250 1570 260
rect 1540 230 1545 250
rect 1565 230 1570 250
rect 1540 200 1570 230
rect 1540 180 1545 200
rect 1565 180 1570 200
rect 1540 170 1570 180
rect 1610 250 1640 260
rect 1610 230 1615 250
rect 1635 230 1640 250
rect 1610 200 1640 230
rect 1610 180 1615 200
rect 1635 180 1640 200
rect 1610 170 1640 180
rect 1665 250 1695 260
rect 1665 230 1670 250
rect 1690 230 1695 250
rect 1665 200 1695 230
rect 1735 250 1765 260
rect 1735 230 1740 250
rect 1760 230 1765 250
rect 1735 200 1765 230
rect 1665 180 1670 200
rect 1690 180 1740 200
rect 1760 180 1765 200
rect 1665 170 1695 180
rect 1735 170 1765 180
rect 1790 250 1820 260
rect 1790 230 1795 250
rect 1815 230 1820 250
rect 1790 200 1820 230
rect 1885 210 1905 300
rect 1940 280 1960 300
rect 1930 275 1970 280
rect 1930 255 1940 275
rect 1960 255 1970 275
rect 1930 250 1970 255
rect 1790 180 1795 200
rect 1815 180 1820 200
rect 1875 205 1970 210
rect 1875 185 1890 205
rect 1910 185 1935 205
rect 1955 185 1970 205
rect 1875 180 1970 185
rect 1790 170 1820 180
rect 1310 140 1350 145
rect 1310 120 1320 140
rect 1340 120 1350 140
rect 1310 115 1350 120
rect 1540 90 1565 170
rect 1615 145 1635 170
rect 1605 140 1645 145
rect 1605 120 1615 140
rect 1635 120 1645 140
rect 1605 115 1645 120
rect 1790 90 1815 170
rect 1355 85 1450 90
rect 1355 65 1370 85
rect 1390 65 1415 85
rect 1435 65 1450 85
rect 1355 60 1450 65
rect 1480 85 1575 90
rect 1480 65 1495 85
rect 1515 65 1540 85
rect 1560 65 1575 85
rect 1480 60 1575 65
rect 1605 85 1700 90
rect 1605 65 1620 85
rect 1640 65 1665 85
rect 1685 65 1700 85
rect 1605 60 1700 65
rect 1730 85 1825 90
rect 1730 65 1745 85
rect 1765 65 1790 85
rect 1810 65 1825 85
rect 1730 60 1825 65
<< viali >>
rect 1415 645 1435 665
rect 1540 645 1560 665
rect 1665 645 1685 665
rect 1790 645 1810 665
rect 1260 585 1280 605
rect 1215 395 1235 415
rect 1935 565 1955 585
rect 1670 380 1690 400
rect 1795 380 1815 400
rect 1890 375 1910 395
rect 1380 335 1400 355
rect 1505 330 1525 350
rect 1265 275 1285 295
rect 1630 290 1650 310
rect 1785 295 1805 315
rect 1260 205 1280 225
rect 1940 255 1960 275
rect 1935 185 1955 205
rect 1320 120 1340 140
rect 1615 120 1635 140
rect 1415 65 1435 85
rect 1540 65 1560 85
rect 1665 65 1685 85
rect 1790 65 1810 85
<< metal1 >>
rect 1115 820 1990 840
rect 1155 700 1195 705
rect 1155 670 1160 700
rect 1190 670 1195 700
rect 1155 665 1195 670
rect 1165 415 1185 665
rect 1260 610 1280 820
rect 1415 670 1435 820
rect 1450 800 1490 805
rect 1450 770 1455 800
rect 1485 770 1490 800
rect 1450 765 1490 770
rect 1405 665 1445 670
rect 1405 645 1415 665
rect 1435 645 1445 665
rect 1405 640 1445 645
rect 1250 605 1290 610
rect 1250 585 1260 605
rect 1280 585 1290 605
rect 1250 580 1290 585
rect 1205 415 1245 420
rect 1165 395 1215 415
rect 1235 395 1325 415
rect 1205 390 1245 395
rect 1305 360 1325 395
rect 1305 355 1410 360
rect 1305 340 1380 355
rect 1370 335 1380 340
rect 1400 335 1410 355
rect 1370 330 1410 335
rect 1460 350 1480 765
rect 1540 670 1560 820
rect 1665 670 1685 820
rect 1790 670 1810 820
rect 1530 665 1570 670
rect 1530 645 1540 665
rect 1560 645 1570 665
rect 1530 640 1570 645
rect 1655 665 1695 670
rect 1655 645 1665 665
rect 1685 645 1695 665
rect 1655 640 1695 645
rect 1780 665 1820 670
rect 1780 645 1790 665
rect 1810 645 1820 665
rect 1780 640 1820 645
rect 1935 590 1955 820
rect 1925 585 1965 590
rect 1925 565 1935 585
rect 1955 565 1965 585
rect 1925 560 1965 565
rect 1660 400 1700 405
rect 1785 400 1825 405
rect 1660 380 1670 400
rect 1690 380 1795 400
rect 1815 395 1825 400
rect 1880 395 1920 400
rect 1815 380 1890 395
rect 1660 375 1700 380
rect 1785 375 1890 380
rect 1910 375 1920 395
rect 1495 350 1535 355
rect 1460 330 1505 350
rect 1525 330 1535 350
rect 1495 325 1535 330
rect 1775 320 1815 325
rect 1570 310 1660 315
rect 1255 295 1295 300
rect 1570 295 1630 310
rect 1255 275 1265 295
rect 1285 275 1590 295
rect 1620 290 1630 295
rect 1650 290 1660 310
rect 1620 285 1660 290
rect 1775 290 1780 320
rect 1810 290 1815 320
rect 1775 285 1815 290
rect 1255 270 1295 275
rect 1250 225 1290 230
rect 1250 205 1260 225
rect 1280 205 1290 225
rect 1250 200 1290 205
rect 1260 -20 1280 200
rect 1310 140 1350 145
rect 1605 140 1645 145
rect 1845 140 1865 375
rect 1880 370 1920 375
rect 1930 275 1970 280
rect 1930 255 1940 275
rect 1960 255 2045 275
rect 1930 250 1970 255
rect 1925 205 1965 210
rect 1925 185 1935 205
rect 1955 185 1965 205
rect 1925 180 1965 185
rect 1310 120 1320 140
rect 1340 120 1615 140
rect 1635 120 1865 140
rect 1310 115 1350 120
rect 1605 115 1645 120
rect 1405 85 1445 90
rect 1405 65 1415 85
rect 1435 65 1445 85
rect 1405 60 1445 65
rect 1530 85 1570 90
rect 1530 65 1540 85
rect 1560 65 1570 85
rect 1530 60 1570 65
rect 1655 85 1695 90
rect 1655 65 1665 85
rect 1685 65 1695 85
rect 1655 60 1695 65
rect 1780 85 1820 90
rect 1780 65 1790 85
rect 1810 65 1820 85
rect 1780 60 1820 65
rect 1415 -20 1435 60
rect 1540 -20 1560 60
rect 1665 -20 1685 60
rect 1790 -20 1810 60
rect 1935 -20 1955 180
rect 1115 -40 1990 -20
<< via1 >>
rect 1160 670 1190 700
rect 1455 770 1485 800
rect 1780 315 1810 320
rect 1780 295 1785 315
rect 1785 295 1805 315
rect 1805 295 1810 315
rect 1780 290 1810 295
<< metal2 >>
rect 1450 800 1490 805
rect 1450 795 1455 800
rect 1115 775 1455 795
rect 1450 770 1455 775
rect 1485 770 1490 800
rect 1450 765 1490 770
rect 1115 725 1725 745
rect 1155 700 1195 705
rect 1155 695 1160 700
rect 1115 675 1160 695
rect 1155 670 1160 675
rect 1190 670 1195 700
rect 1155 665 1195 670
rect 1705 305 1725 725
rect 1775 320 1815 325
rect 1775 305 1780 320
rect 1705 290 1780 305
rect 1810 290 1815 320
rect 1705 285 1815 290
<< labels >>
rlabel metal2 1120 675 1130 695 1 sel
rlabel metal2 1120 725 1130 745 1 in1
rlabel metal2 1120 775 1130 795 1 in2
rlabel metal1 1240 830 1240 830 1 vdd
rlabel metal1 2030 255 2040 275 1 out
rlabel metal1 1235 -30 1235 -30 1 gnd
<< end >>
