magic
tech sky130A
timestamp 1720964864
<< metal1 >>
rect 2015 935 4610 955
rect 2195 900 2235 905
rect 2195 870 2200 900
rect 2230 870 2235 900
rect 2195 865 2235 870
rect 4485 900 4525 905
rect 4485 870 4490 900
rect 4520 870 4525 900
rect 4485 865 4525 870
rect 6775 900 6815 905
rect 6775 870 6780 900
rect 6810 870 6815 900
rect 6775 865 6815 870
rect 2090 420 2130 425
rect 2090 390 2095 420
rect 2125 390 2130 420
rect 2090 385 2130 390
rect 2205 365 2225 865
rect 4380 420 4420 425
rect 4310 385 4330 400
rect 4380 390 4385 420
rect 4415 390 4420 420
rect 4380 385 4420 390
rect 4495 365 4515 865
rect 6670 420 6710 425
rect 6670 405 6675 420
rect 6650 390 6675 405
rect 6705 390 6710 420
rect 6650 385 6710 390
rect 6785 365 6805 865
rect 8960 420 9000 425
rect 8960 390 8965 420
rect 8995 390 9000 420
rect 8960 385 9000 390
rect 2090 345 2225 365
rect 4380 345 4515 365
rect 6665 345 6805 365
rect 2015 0 6885 20
rect -540 -45 -500 -40
rect -540 -75 -535 -45
rect -505 -75 -500 -45
rect -540 -80 -500 -75
rect -530 -1330 -510 -80
rect -480 -95 -440 -90
rect -480 -125 -475 -95
rect -445 -125 -440 -95
rect -480 -130 -440 -125
rect -540 -1335 -500 -1330
rect -540 -1365 -535 -1335
rect -505 -1365 -500 -1335
rect -540 -1370 -500 -1365
rect -470 -1380 -450 -130
rect -420 -145 -380 -140
rect -420 -175 -415 -145
rect -385 -175 -380 -145
rect -420 -180 -380 -175
rect -480 -1385 -440 -1380
rect -480 -1415 -475 -1385
rect -445 -1415 -440 -1385
rect -480 -1420 -440 -1415
rect -410 -1430 -390 -180
rect -360 -195 -320 -190
rect -360 -225 -355 -195
rect -325 -225 -320 -195
rect -360 -230 -320 -225
rect -420 -1435 -380 -1430
rect -420 -1465 -415 -1435
rect -385 -1465 -380 -1435
rect -420 -1470 -380 -1465
rect -350 -1480 -330 -230
rect -300 -245 -260 -240
rect -300 -275 -295 -245
rect -265 -275 -260 -245
rect -300 -280 -260 -275
rect -360 -1485 -320 -1480
rect -360 -1515 -355 -1485
rect -325 -1515 -320 -1485
rect -360 -1520 -320 -1515
rect -290 -1530 -270 -280
rect -240 -295 -200 -290
rect -240 -325 -235 -295
rect -205 -325 -200 -295
rect -240 -330 -200 -325
rect -300 -1535 -260 -1530
rect -300 -1565 -295 -1535
rect -265 -1565 -260 -1535
rect -300 -1570 -260 -1565
rect -230 -1580 -210 -330
rect 1760 -340 1835 -335
rect 1895 -340 2000 -335
rect 2015 -355 6875 -335
rect 2195 -390 2235 -385
rect 2195 -420 2200 -390
rect 2230 -420 2235 -390
rect 2195 -425 2235 -420
rect 4485 -390 4525 -385
rect 4485 -420 4490 -390
rect 4520 -420 4525 -390
rect 4485 -425 4525 -420
rect 6775 -390 6815 -385
rect 6775 -420 6780 -390
rect 6810 -420 6815 -390
rect 6775 -425 6815 -420
rect -120 -440 -80 -435
rect -120 -470 -115 -440
rect -85 -470 -80 -440
rect -120 -475 -80 -470
rect -180 -540 -140 -535
rect -180 -570 -175 -540
rect -145 -570 -140 -540
rect -180 -575 -140 -570
rect -240 -1585 -200 -1580
rect -240 -1615 -235 -1585
rect -205 -1615 -200 -1585
rect -240 -1620 -200 -1615
rect -170 -1675 -150 -575
rect -180 -1680 -140 -1675
rect -180 -1710 -175 -1680
rect -145 -1710 -140 -1680
rect -180 -1715 -140 -1710
rect -110 -1725 -90 -475
rect -60 -490 -20 -485
rect -60 -520 -55 -490
rect -25 -520 -20 -490
rect -60 -525 -20 -520
rect -120 -1730 -80 -1725
rect -120 -1760 -115 -1730
rect -85 -1760 -80 -1730
rect -120 -1765 -80 -1760
rect -50 -1775 -30 -525
rect 2090 -870 2130 -865
rect 2090 -900 2095 -870
rect 2125 -900 2130 -870
rect 2090 -905 2130 -900
rect 2205 -925 2225 -425
rect 4380 -870 4420 -865
rect 4380 -900 4385 -870
rect 4415 -900 4420 -870
rect 4380 -905 4420 -900
rect 4495 -925 4515 -425
rect 6670 -870 6710 -865
rect 6670 -900 6675 -870
rect 6705 -900 6710 -870
rect 6670 -905 6710 -900
rect 6785 -925 6805 -425
rect 8945 -830 8960 365
rect 8945 -845 9135 -830
rect 8960 -870 9000 -865
rect 8960 -900 8965 -870
rect 8995 -900 9000 -870
rect 8960 -905 9000 -900
rect 9065 -920 9105 -915
rect 9065 -925 9070 -920
rect 2090 -945 2225 -925
rect 4380 -945 4515 -925
rect 6670 -945 6805 -925
rect 8960 -945 9070 -925
rect 9065 -950 9070 -945
rect 9100 -950 9105 -920
rect 9065 -955 9105 -950
rect 2015 -1290 6870 -1270
rect 2090 -1330 2130 -1325
rect 2090 -1360 2095 -1330
rect 2125 -1360 2130 -1330
rect 2090 -1365 2130 -1360
rect 4380 -1330 4420 -1325
rect 4380 -1360 4385 -1330
rect 4415 -1360 4420 -1330
rect 4380 -1365 4420 -1360
rect 6670 -1330 6710 -1325
rect 6670 -1360 6675 -1330
rect 6705 -1360 6710 -1330
rect 6670 -1365 6710 -1360
rect 8960 -1330 9000 -1325
rect 8960 -1360 8965 -1330
rect 8995 -1360 9000 -1330
rect 8960 -1365 9000 -1360
rect 2100 -1625 2120 -1365
rect 4390 -1625 4410 -1365
rect 6680 -1625 6700 -1365
rect 1780 -1630 1835 -1625
rect 1940 -1630 6880 -1625
rect 2005 -1645 6880 -1630
rect -60 -1780 -20 -1775
rect -60 -1810 -55 -1780
rect -25 -1810 -20 -1780
rect -60 -1815 -20 -1810
rect 2100 -1945 2120 -1645
rect 2195 -1680 2235 -1675
rect 2195 -1710 2200 -1680
rect 2230 -1710 2235 -1680
rect 2195 -1715 2235 -1710
rect 2090 -1950 2130 -1945
rect 2090 -1980 2095 -1950
rect 2125 -1980 2130 -1950
rect 2090 -1985 2130 -1980
rect 2150 -2160 2190 -2155
rect 2150 -2175 2155 -2160
rect 2090 -2190 2155 -2175
rect 2185 -2190 2190 -2160
rect 2090 -2195 2190 -2190
rect 2205 -2215 2225 -1715
rect 4390 -1945 4410 -1645
rect 4485 -1680 4525 -1675
rect 4485 -1710 4490 -1680
rect 4520 -1710 4525 -1680
rect 4485 -1715 4525 -1710
rect 4380 -1950 4420 -1945
rect 4380 -1980 4385 -1950
rect 4415 -1980 4420 -1950
rect 4380 -1985 4420 -1980
rect 4440 -2160 4480 -2155
rect 4440 -2175 4445 -2160
rect 4380 -2190 4445 -2175
rect 4475 -2190 4480 -2160
rect 4380 -2195 4480 -2190
rect 4495 -2215 4515 -1715
rect 6680 -1945 6700 -1645
rect 6775 -1680 6815 -1675
rect 6775 -1710 6780 -1680
rect 6810 -1710 6815 -1680
rect 6775 -1715 6815 -1710
rect 6670 -1950 6710 -1945
rect 6670 -1980 6675 -1950
rect 6705 -1980 6710 -1950
rect 6670 -1985 6710 -1980
rect 6730 -2160 6770 -2155
rect 6730 -2175 6735 -2160
rect 6670 -2190 6735 -2175
rect 6765 -2190 6770 -2160
rect 6670 -2195 6770 -2190
rect 6785 -2215 6805 -1715
rect 8970 -1945 8990 -1365
rect 8960 -1950 9000 -1945
rect 8960 -1980 8965 -1950
rect 8995 -1980 9000 -1950
rect 8960 -1985 9000 -1980
rect 9020 -2160 9060 -2155
rect 9020 -2175 9025 -2160
rect 8960 -2190 9025 -2175
rect 9055 -2190 9060 -2160
rect 9120 -2170 9135 -845
rect 9120 -2185 9175 -2170
rect 8960 -2195 9060 -2190
rect 9105 -2210 9145 -2205
rect 9105 -2215 9110 -2210
rect 2090 -2235 2225 -2215
rect 4380 -2235 4515 -2215
rect 6670 -2235 6805 -2215
rect 8950 -2235 9110 -2215
rect 9105 -2240 9110 -2235
rect 9140 -2240 9145 -2210
rect 9105 -2245 9145 -2240
rect 9160 -2275 9175 -2185
rect 9030 -2290 9175 -2275
rect 2015 -2580 6885 -2560
rect 870 -2885 8125 -2865
rect 9030 -2900 9050 -2290
rect 9020 -2905 9060 -2900
rect 9020 -2935 9025 -2905
rect 9055 -2935 9060 -2905
rect 9020 -2940 9060 -2935
rect 910 -3660 930 -3430
rect 2845 -3450 2920 -3430
rect 4835 -3450 4910 -3430
rect 6825 -3450 6900 -3430
rect 8815 -3450 8890 -3430
rect 2900 -3660 2920 -3450
rect 4890 -3660 4910 -3450
rect 6880 -3660 6900 -3450
rect 8870 -3660 8890 -3450
rect 900 -3665 940 -3660
rect 900 -3695 905 -3665
rect 935 -3695 940 -3665
rect 900 -3700 940 -3695
rect 2890 -3665 2930 -3660
rect 2890 -3695 2895 -3665
rect 2925 -3695 2930 -3665
rect 2890 -3700 2930 -3695
rect 4880 -3665 4920 -3660
rect 4880 -3695 4885 -3665
rect 4915 -3695 4920 -3665
rect 4880 -3700 4920 -3695
rect 6870 -3665 6910 -3660
rect 6870 -3695 6875 -3665
rect 6905 -3695 6910 -3665
rect 6870 -3700 6910 -3695
rect 8860 -3665 8900 -3660
rect 8860 -3695 8865 -3665
rect 8895 -3695 8900 -3665
rect 8860 -3700 8900 -3695
rect 875 -3745 7975 -3725
<< via1 >>
rect 2200 870 2230 900
rect 4490 870 4520 900
rect 6780 870 6810 900
rect 2095 390 2125 420
rect 4385 390 4415 420
rect 6675 390 6705 420
rect 8965 390 8995 420
rect -535 -75 -505 -45
rect -475 -125 -445 -95
rect -535 -1365 -505 -1335
rect -415 -175 -385 -145
rect -475 -1415 -445 -1385
rect -355 -225 -325 -195
rect -415 -1465 -385 -1435
rect -295 -275 -265 -245
rect -355 -1515 -325 -1485
rect -235 -325 -205 -295
rect -295 -1565 -265 -1535
rect 2200 -420 2230 -390
rect 4490 -420 4520 -390
rect 6780 -420 6810 -390
rect -115 -470 -85 -440
rect -175 -570 -145 -540
rect -235 -1615 -205 -1585
rect -175 -1710 -145 -1680
rect -55 -520 -25 -490
rect -115 -1760 -85 -1730
rect 2095 -900 2125 -870
rect 4385 -900 4415 -870
rect 6675 -900 6705 -870
rect 8965 -900 8995 -870
rect 9070 -950 9100 -920
rect 2095 -1360 2125 -1330
rect 4385 -1360 4415 -1330
rect 6675 -1360 6705 -1330
rect 8965 -1360 8995 -1330
rect -55 -1810 -25 -1780
rect 2200 -1710 2230 -1680
rect 2095 -1980 2125 -1950
rect 2155 -2190 2185 -2160
rect 4490 -1710 4520 -1680
rect 4385 -1980 4415 -1950
rect 4445 -2190 4475 -2160
rect 6780 -1710 6810 -1680
rect 6675 -1980 6705 -1950
rect 6735 -2190 6765 -2160
rect 8965 -1980 8995 -1950
rect 9025 -2190 9055 -2160
rect 9110 -2240 9140 -2210
rect 9025 -2935 9055 -2905
rect 905 -3695 935 -3665
rect 2895 -3695 2925 -3665
rect 4885 -3695 4915 -3665
rect 6875 -3695 6905 -3665
rect 8865 -3695 8895 -3665
<< metal2 >>
rect -620 1130 6710 1150
rect -620 1095 6670 1115
rect -620 1060 4420 1080
rect -620 1025 4380 1045
rect -620 990 2130 1010
rect -620 955 2090 975
rect 2110 955 2130 990
rect 4360 955 4380 1025
rect 4400 955 4420 1060
rect -620 920 5 940
rect -620 885 -35 905
rect -620 850 -75 870
rect -95 795 -75 850
rect -55 845 -35 885
rect -15 875 5 920
rect -55 825 5 845
rect 2070 795 2090 935
rect 2110 845 2130 935
rect 2195 900 2235 905
rect 2195 870 2200 900
rect 2230 895 2235 900
rect 2230 875 2295 895
rect 2230 870 2235 875
rect 2195 865 2235 870
rect 2110 825 2295 845
rect 4360 795 4380 935
rect 4400 845 4420 935
rect 4485 900 4525 905
rect 4485 870 4490 900
rect 4520 895 4525 900
rect 4520 875 4585 895
rect 4520 870 4525 875
rect 4485 865 4525 870
rect 4400 825 4585 845
rect 6650 795 6670 1095
rect 6690 845 6710 1130
rect 6775 900 6815 905
rect 6775 870 6780 900
rect 6810 895 6815 900
rect 6810 875 6875 895
rect 6810 870 6815 875
rect 6775 865 6815 870
rect 6690 825 6875 845
rect -95 775 5 795
rect 2070 775 2295 795
rect 4360 775 4585 795
rect 6650 775 6880 795
rect 2090 420 2130 425
rect 2090 390 2095 420
rect 2125 390 2130 420
rect 2090 385 2130 390
rect 4380 420 4420 425
rect 4380 390 4385 420
rect 4415 390 4420 420
rect 4380 385 4420 390
rect 6670 420 6710 425
rect 6670 390 6675 420
rect 6705 390 6710 420
rect 6670 385 6710 390
rect 8960 420 9000 425
rect 8960 390 8965 420
rect 8995 390 9000 420
rect 8960 385 9000 390
rect -540 -45 -500 -40
rect -540 -50 -535 -45
rect -625 -70 -535 -50
rect -540 -75 -535 -70
rect -505 -50 -500 -45
rect -505 -70 1830 -50
rect -505 -75 -500 -70
rect -540 -80 -500 -75
rect -480 -95 -440 -90
rect -480 -100 -475 -95
rect -625 -120 -475 -100
rect -480 -125 -475 -120
rect -445 -100 -440 -95
rect -445 -120 1790 -100
rect -445 -125 -440 -120
rect -480 -130 -440 -125
rect -420 -145 -380 -140
rect -420 -150 -415 -145
rect -625 -170 -415 -150
rect -420 -175 -415 -170
rect -385 -150 -380 -145
rect -385 -170 1750 -150
rect -385 -175 -380 -170
rect -420 -180 -380 -175
rect -360 -195 -320 -190
rect -360 -200 -355 -195
rect -625 -220 -355 -200
rect -360 -225 -355 -220
rect -325 -200 -320 -195
rect -325 -220 1710 -200
rect -325 -225 -320 -220
rect -360 -230 -320 -225
rect -300 -245 -260 -240
rect -300 -250 -295 -245
rect -625 -270 -295 -250
rect -300 -275 -295 -270
rect -265 -250 -260 -245
rect 1690 -245 1710 -220
rect 1730 -210 1750 -170
rect 1770 -175 1790 -120
rect 1810 -140 1830 -70
rect 2100 -105 2120 385
rect 4390 -70 4410 385
rect 6680 -35 6700 385
rect 8970 0 8990 385
rect 8970 -20 9090 0
rect 6680 -55 9090 -35
rect 4390 -90 9090 -70
rect 2100 -125 9090 -105
rect 1810 -160 6710 -140
rect 1770 -195 6670 -175
rect 1730 -230 4420 -210
rect -265 -270 1670 -250
rect 1690 -265 4380 -245
rect -265 -275 -260 -270
rect -300 -280 -260 -275
rect 1650 -280 1670 -270
rect -240 -295 -200 -290
rect -240 -300 -235 -295
rect -625 -320 -235 -300
rect -240 -325 -235 -320
rect -205 -300 -200 -295
rect 1650 -300 2130 -280
rect -205 -315 1630 -300
rect -205 -320 2090 -315
rect -205 -325 -200 -320
rect -240 -330 -200 -325
rect 1610 -335 2090 -320
rect -625 -415 5 -395
rect -120 -440 -80 -435
rect -120 -445 -115 -440
rect -625 -465 -115 -445
rect -120 -470 -115 -465
rect -85 -445 -80 -440
rect -85 -465 5 -445
rect -85 -470 -80 -465
rect -120 -475 -80 -470
rect -60 -490 -20 -485
rect -60 -495 -55 -490
rect -625 -515 -55 -495
rect -60 -520 -55 -515
rect -25 -495 -20 -490
rect 2070 -495 2090 -335
rect 2110 -445 2130 -300
rect 2195 -390 2235 -385
rect 2195 -420 2200 -390
rect 2230 -395 2235 -390
rect 2230 -415 2295 -395
rect 2230 -420 2235 -415
rect 2195 -425 2235 -420
rect 2110 -465 2295 -445
rect 4360 -495 4380 -265
rect 4400 -445 4420 -230
rect 4485 -390 4525 -385
rect 4485 -420 4490 -390
rect 4520 -395 4525 -390
rect 4520 -415 4585 -395
rect 4520 -420 4525 -415
rect 4485 -425 4525 -420
rect 4400 -465 4585 -445
rect 6650 -495 6670 -195
rect 6690 -445 6710 -160
rect 6775 -390 6815 -385
rect 6775 -420 6780 -390
rect 6810 -395 6815 -390
rect 6810 -415 6875 -395
rect 6810 -420 6815 -415
rect 6775 -425 6815 -420
rect 6690 -465 6875 -445
rect -25 -515 5 -495
rect 2070 -515 2295 -495
rect 4360 -515 4585 -495
rect 6650 -515 6875 -495
rect -25 -520 -20 -515
rect -60 -525 -20 -520
rect -180 -540 -140 -535
rect -180 -545 -175 -540
rect -625 -565 -175 -545
rect -180 -570 -175 -565
rect -145 -570 -140 -540
rect -180 -575 -140 -570
rect 2090 -870 2130 -865
rect 2090 -900 2095 -870
rect 2125 -900 2130 -870
rect 2090 -905 2130 -900
rect 4380 -870 4420 -865
rect 4380 -900 4385 -870
rect 4415 -900 4420 -870
rect 4380 -905 4420 -900
rect 6670 -870 6710 -865
rect 6670 -900 6675 -870
rect 6705 -900 6710 -870
rect 6670 -905 6710 -900
rect 8960 -870 9000 -865
rect 8960 -900 8965 -870
rect 8995 -900 9000 -870
rect 8960 -905 9000 -900
rect 2100 -1325 2120 -905
rect 4390 -1325 4410 -905
rect 6680 -1325 6700 -905
rect 8970 -1325 8990 -905
rect 9065 -920 9105 -915
rect 9065 -950 9070 -920
rect 9100 -950 9105 -920
rect 9065 -955 9105 -950
rect 2090 -1330 2130 -1325
rect -540 -1335 -500 -1330
rect -540 -1365 -535 -1335
rect -505 -1340 -500 -1335
rect -505 -1360 1830 -1340
rect -505 -1365 -500 -1360
rect -540 -1370 -500 -1365
rect -480 -1385 -440 -1380
rect -480 -1415 -475 -1385
rect -445 -1390 -440 -1385
rect -445 -1410 1790 -1390
rect -445 -1415 -440 -1410
rect -480 -1420 -440 -1415
rect -420 -1435 -380 -1430
rect -420 -1465 -415 -1435
rect -385 -1440 -380 -1435
rect -385 -1460 1750 -1440
rect -385 -1465 -380 -1460
rect -420 -1470 -380 -1465
rect -360 -1485 -320 -1480
rect -360 -1515 -355 -1485
rect -325 -1490 -320 -1485
rect -325 -1510 1710 -1490
rect -325 -1515 -320 -1510
rect -360 -1520 -320 -1515
rect -300 -1535 -260 -1530
rect -300 -1565 -295 -1535
rect -265 -1540 -260 -1535
rect 1690 -1535 1710 -1510
rect 1730 -1500 1750 -1460
rect 1770 -1465 1790 -1410
rect 1810 -1430 1830 -1360
rect 2090 -1360 2095 -1330
rect 2125 -1360 2130 -1330
rect 2090 -1365 2130 -1360
rect 4380 -1330 4420 -1325
rect 4380 -1360 4385 -1330
rect 4415 -1360 4420 -1330
rect 4380 -1365 4420 -1360
rect 6670 -1330 6710 -1325
rect 6670 -1360 6675 -1330
rect 6705 -1360 6710 -1330
rect 6670 -1365 6710 -1360
rect 8960 -1330 9000 -1325
rect 8960 -1360 8965 -1330
rect 8995 -1360 9000 -1330
rect 8960 -1365 9000 -1360
rect 1810 -1450 6710 -1430
rect 1770 -1485 6670 -1465
rect 1730 -1520 4420 -1500
rect -265 -1560 1670 -1540
rect 1690 -1555 4380 -1535
rect -265 -1565 -260 -1560
rect -300 -1570 -260 -1565
rect 1650 -1570 1670 -1560
rect -240 -1585 -200 -1580
rect -240 -1615 -235 -1585
rect -205 -1590 -200 -1585
rect 1650 -1590 2130 -1570
rect -205 -1605 1630 -1590
rect -205 -1610 2090 -1605
rect -205 -1615 -200 -1610
rect -240 -1620 -200 -1615
rect 1610 -1625 2090 -1610
rect -180 -1680 -140 -1675
rect -180 -1710 -175 -1680
rect -145 -1685 -140 -1680
rect -145 -1705 5 -1685
rect -145 -1710 -140 -1705
rect -180 -1715 -140 -1710
rect -120 -1730 -80 -1725
rect -120 -1760 -115 -1730
rect -85 -1735 -80 -1730
rect -85 -1755 5 -1735
rect -85 -1760 -80 -1755
rect -120 -1765 -80 -1760
rect -60 -1780 -20 -1775
rect -60 -1810 -55 -1780
rect -25 -1785 -20 -1780
rect 2070 -1785 2090 -1625
rect 2110 -1735 2130 -1590
rect 2195 -1680 2235 -1675
rect 2195 -1710 2200 -1680
rect 2230 -1685 2235 -1680
rect 2230 -1705 2295 -1685
rect 2230 -1710 2235 -1705
rect 2195 -1715 2235 -1710
rect 2110 -1755 2295 -1735
rect 4360 -1785 4380 -1555
rect 4400 -1735 4420 -1520
rect 4485 -1680 4525 -1675
rect 4485 -1710 4490 -1680
rect 4520 -1685 4525 -1680
rect 4520 -1705 4585 -1685
rect 4520 -1710 4525 -1705
rect 4485 -1715 4525 -1710
rect 4400 -1755 4585 -1735
rect 6650 -1785 6670 -1485
rect 6690 -1735 6710 -1450
rect 6775 -1680 6815 -1675
rect 6775 -1710 6780 -1680
rect 6810 -1685 6815 -1680
rect 6810 -1705 6875 -1685
rect 6810 -1710 6815 -1705
rect 6775 -1715 6815 -1710
rect 6690 -1755 6875 -1735
rect -25 -1805 5 -1785
rect 2070 -1805 2295 -1785
rect 4360 -1805 4585 -1785
rect 6650 -1805 6875 -1785
rect -25 -1810 -20 -1805
rect -60 -1815 -20 -1810
rect 2090 -1950 2130 -1945
rect 2090 -1980 2095 -1950
rect 2125 -1980 2130 -1950
rect 2090 -1985 2130 -1980
rect 4380 -1950 4420 -1945
rect 4380 -1980 4385 -1950
rect 4415 -1980 4420 -1950
rect 4380 -1985 4420 -1980
rect 6670 -1950 6710 -1945
rect 6670 -1980 6675 -1950
rect 6705 -1980 6710 -1950
rect 6670 -1985 6710 -1980
rect 8960 -1950 9000 -1945
rect 8960 -1980 8965 -1950
rect 8995 -1980 9000 -1950
rect 8960 -1985 9000 -1980
rect 2100 -2580 2120 -1985
rect 2150 -2160 2190 -2155
rect 2150 -2190 2155 -2160
rect 2185 -2190 2190 -2160
rect 2150 -2195 2190 -2190
rect -80 -2595 2120 -2580
rect -80 -2960 -60 -2595
rect 2160 -2610 2180 -2195
rect -45 -2625 2180 -2610
rect -45 -2910 -25 -2625
rect 4390 -2640 4410 -1985
rect 4440 -2160 4480 -2155
rect 4440 -2190 4445 -2160
rect 4475 -2190 4480 -2160
rect 4440 -2195 4480 -2190
rect 1910 -2655 4410 -2640
rect -45 -2930 0 -2910
rect 1910 -2960 1930 -2655
rect 4450 -2670 4470 -2195
rect 1945 -2685 4470 -2670
rect 1945 -2910 1965 -2685
rect 6680 -2700 6700 -1985
rect 6730 -2160 6770 -2155
rect 6730 -2190 6735 -2160
rect 6765 -2190 6770 -2160
rect 6730 -2195 6770 -2190
rect 3900 -2715 6700 -2700
rect 1945 -2930 1990 -2910
rect 3900 -2960 3920 -2715
rect 6740 -2730 6760 -2195
rect 3935 -2745 6760 -2730
rect 3935 -2910 3955 -2745
rect 8970 -2760 8990 -1985
rect 9020 -2160 9060 -2155
rect 9020 -2190 9025 -2160
rect 9055 -2190 9060 -2160
rect 9020 -2195 9060 -2190
rect 5890 -2775 8990 -2760
rect 3935 -2930 3980 -2910
rect 5890 -2960 5910 -2775
rect 9030 -2790 9050 -2195
rect 5925 -2805 9050 -2790
rect 5925 -2910 5945 -2805
rect 9075 -2820 9090 -955
rect 9105 -2210 9145 -2205
rect 9105 -2240 9110 -2210
rect 9140 -2240 9145 -2210
rect 9105 -2245 9145 -2240
rect 7885 -2835 9090 -2820
rect 5925 -2930 5970 -2910
rect 7885 -2960 7905 -2835
rect 9115 -2850 9135 -2245
rect 7920 -2865 9135 -2850
rect 7920 -2910 7940 -2865
rect 9020 -2905 9060 -2900
rect 7920 -2930 7965 -2910
rect 9020 -2935 9025 -2905
rect 9055 -2935 9060 -2905
rect 9020 -2940 9060 -2935
rect -80 -2980 0 -2960
rect 1910 -2980 1990 -2960
rect 3900 -2980 3980 -2960
rect 5890 -2980 5970 -2960
rect 7885 -2980 7965 -2960
rect -80 -3030 0 -3010
rect 1910 -3030 1990 -3010
rect 3900 -3030 3980 -3010
rect 5890 -3030 5970 -3010
rect 7885 -3030 7960 -3010
rect -80 -3630 -60 -3030
rect 1910 -3630 1930 -3030
rect 3900 -3630 3920 -3030
rect 5890 -3630 5910 -3030
rect 7885 -3630 7900 -3030
rect 9030 -3630 9050 -2940
rect -80 -3645 9050 -3630
rect 900 -3665 940 -3660
rect 900 -3695 905 -3665
rect 935 -3695 940 -3665
rect 900 -3700 940 -3695
rect 2890 -3665 2930 -3660
rect 2890 -3695 2895 -3665
rect 2925 -3695 2930 -3665
rect 2890 -3700 2930 -3695
rect 4880 -3665 4920 -3660
rect 4880 -3695 4885 -3665
rect 4915 -3695 4920 -3665
rect 4880 -3700 4920 -3695
rect 6870 -3665 6910 -3660
rect 6870 -3695 6875 -3665
rect 6905 -3695 6910 -3665
rect 6870 -3700 6910 -3695
rect 8860 -3665 8900 -3660
rect 8860 -3695 8865 -3665
rect 8895 -3670 8900 -3665
rect 8895 -3690 9140 -3670
rect 8895 -3695 8900 -3690
rect 8860 -3700 8900 -3695
rect 910 -3820 930 -3700
rect 2900 -3785 2920 -3700
rect 4890 -3750 4910 -3700
rect 6880 -3715 6900 -3700
rect 6880 -3735 9140 -3715
rect 4890 -3770 9140 -3750
rect 2900 -3805 9140 -3785
rect 910 -3840 9140 -3820
use full_adder  full_adder_0
timestamp 1720949016
transform 1 0 2380 0 1 460
box -90 -460 2000 495
use full_adder  full_adder_1
timestamp 1720949016
transform 1 0 90 0 1 460
box -90 -460 2000 495
use full_adder  full_adder_2
timestamp 1720949016
transform 1 0 4670 0 1 460
box -90 -460 2000 495
use full_adder  full_adder_3
timestamp 1720949016
transform 1 0 6960 0 1 -830
box -90 -460 2000 495
use full_adder  full_adder_4
timestamp 1720949016
transform 1 0 6960 0 1 460
box -90 -460 2000 495
use full_adder  full_adder_5
timestamp 1720949016
transform 1 0 90 0 1 -830
box -90 -460 2000 495
use full_adder  full_adder_6
timestamp 1720949016
transform 1 0 2380 0 1 -830
box -90 -460 2000 495
use full_adder  full_adder_7
timestamp 1720949016
transform 1 0 4670 0 1 -830
box -90 -460 2000 495
use full_adder  full_adder_8
timestamp 1720949016
transform 1 0 2380 0 1 -2120
box -90 -460 2000 495
use full_adder  full_adder_9
timestamp 1720949016
transform 1 0 90 0 1 -2120
box -90 -460 2000 495
use full_adder  full_adder_10
timestamp 1720949016
transform 1 0 4670 0 1 -2120
box -90 -460 2000 495
use full_adder  full_adder_11
timestamp 1720949016
transform 1 0 6960 0 1 -2120
box -90 -460 2000 495
use mux_2to1  mux_2to1_0
timestamp 1720937323
transform 1 0 -1115 0 1 -3705
box 1115 -40 2045 840
use mux_2to1  mux_2to1_1
timestamp 1720937323
transform 1 0 875 0 1 -3705
box 1115 -40 2045 840
use mux_2to1  mux_2to1_2
timestamp 1720937323
transform 1 0 2865 0 1 -3705
box 1115 -40 2045 840
use mux_2to1  mux_2to1_3
timestamp 1720937323
transform 1 0 4855 0 1 -3705
box 1115 -40 2045 840
use mux_2to1  mux_2to1_4
timestamp 1720937323
transform 1 0 6845 0 1 -3705
box 1115 -40 2045 840
<< labels >>
rlabel metal2 -610 850 -600 870 1 a0
rlabel metal2 -610 885 -600 905 1 b0
rlabel metal2 -610 955 -600 975 1 a1
rlabel metal2 -610 1025 -600 1045 1 a2
rlabel metal2 -610 1095 -600 1115 1 a3
rlabel metal2 -610 990 -600 1010 1 b1
rlabel metal2 -610 1060 -600 1080 1 b2
rlabel metal2 -610 1130 -600 1150 1 b3
rlabel metal2 -615 -415 -605 -395 1 cin0
rlabel metal2 -615 -515 -605 -495 1 a4
rlabel metal2 -615 -320 -605 -300 1 a5
rlabel metal2 -615 -220 -605 -200 1 a6
rlabel metal2 -615 -120 -605 -100 1 a7
rlabel metal2 -615 -465 -605 -445 1 b4
rlabel metal2 -615 -270 -605 -250 1 b5
rlabel metal2 -615 -170 -605 -150 1 b6
rlabel metal2 -615 -70 -605 -50 1 b7
rlabel metal2 -615 -565 -605 -545 1 cin1
rlabel metal2 -610 920 -600 940 1 cin0
rlabel metal1 2905 -3450 2915 -3430 1 out
rlabel metal1 4895 -3450 4905 -3430 1 out
rlabel metal1 6885 -3450 6895 -3430 1 out
rlabel metal1 8875 -3450 8885 -3430 1 out
rlabel metal2 9125 -3690 9135 -3670 1 cout
rlabel metal2 9125 -3735 9135 -3715 1 s7
rlabel metal2 9125 -3770 9135 -3750 1 s6
rlabel metal2 9125 -3805 9135 -3785 1 s5
rlabel metal2 9125 -3840 9135 -3820 1 s4
rlabel metal1 6825 -1285 6825 -1285 1 gnd
rlabel metal1 6775 -345 6775 -345 1 vdd
rlabel metal1 6765 5 6765 5 1 gnd
rlabel metal1 4550 945 4550 945 1 vdd
rlabel metal1 2170 -1635 2170 -1635 1 vdd
rlabel metal1 6730 -2575 6730 -2575 1 gnd
rlabel metal1 7800 -2880 7800 -2880 1 vdd
rlabel metal1 7680 -3740 7680 -3740 1 gnd
rlabel metal2 9075 -20 9085 0 1 s3
rlabel metal2 9075 -55 9085 -35 1 s2
rlabel metal2 9075 -90 9085 -70 1 s1
rlabel metal2 9075 -125 9085 -105 1 s0
<< end >>
