magic
tech sky130A
timestamp 1720529296
<< metal1 >>
rect 1775 935 1960 955
rect 3730 935 3905 955
rect 5680 935 5855 955
rect 1915 900 1955 905
rect 1915 870 1920 900
rect 1950 870 1955 900
rect 1915 865 1955 870
rect 3865 900 3905 905
rect 3865 870 3870 900
rect 3900 870 3905 900
rect 3865 865 3905 870
rect 5815 900 5855 905
rect 5815 870 5820 900
rect 5850 870 5855 900
rect 5815 865 5855 870
rect 1855 420 1895 425
rect 1855 390 1860 420
rect 1890 390 1895 420
rect 1855 385 1895 390
rect 1925 365 1945 865
rect 3805 420 3845 425
rect 3805 390 3810 420
rect 3840 390 3845 420
rect 3805 385 3845 390
rect 3875 365 3895 865
rect 5755 420 5795 425
rect 5755 390 5760 420
rect 5790 390 5795 420
rect 5755 385 5795 390
rect 5825 365 5845 865
rect 7705 420 7745 425
rect 7705 390 7710 420
rect 7740 390 7745 420
rect 7705 385 7745 390
rect 1895 345 1945 365
rect 3845 345 3895 365
rect 5795 345 5845 365
rect 7745 345 8000 365
rect 1775 0 5855 20
rect -540 -45 -500 -40
rect -540 -75 -535 -45
rect -505 -75 -500 -45
rect -540 -80 -500 -75
rect -530 -1330 -510 -80
rect -480 -95 -440 -90
rect -480 -125 -475 -95
rect -445 -125 -440 -95
rect -480 -130 -440 -125
rect -540 -1335 -500 -1330
rect -540 -1365 -535 -1335
rect -505 -1365 -500 -1335
rect -540 -1370 -500 -1365
rect -470 -1380 -450 -130
rect -420 -145 -380 -140
rect -420 -175 -415 -145
rect -385 -175 -380 -145
rect -420 -180 -380 -175
rect -480 -1385 -440 -1380
rect -480 -1415 -475 -1385
rect -445 -1415 -440 -1385
rect -480 -1420 -440 -1415
rect -410 -1430 -390 -180
rect -360 -195 -320 -190
rect -360 -225 -355 -195
rect -325 -225 -320 -195
rect -360 -230 -320 -225
rect -420 -1435 -380 -1430
rect -420 -1465 -415 -1435
rect -385 -1465 -380 -1435
rect -420 -1470 -380 -1465
rect -350 -1480 -330 -230
rect -300 -245 -260 -240
rect -300 -275 -295 -245
rect -265 -275 -260 -245
rect -300 -280 -260 -275
rect -360 -1485 -320 -1480
rect -360 -1515 -355 -1485
rect -325 -1515 -320 -1485
rect -360 -1520 -320 -1515
rect -290 -1530 -270 -280
rect -240 -295 -200 -290
rect -240 -325 -235 -295
rect -205 -325 -200 -295
rect -240 -330 -200 -325
rect -300 -1535 -260 -1530
rect -300 -1565 -295 -1535
rect -265 -1565 -260 -1535
rect -300 -1570 -260 -1565
rect -230 -1580 -210 -330
rect 1760 -355 3925 -335
rect 1945 -390 1985 -385
rect 1945 -420 1950 -390
rect 1980 -420 1985 -390
rect 1945 -425 1985 -420
rect 3900 -390 3940 -385
rect 3900 -420 3905 -390
rect 3935 -420 3940 -390
rect 3900 -425 3940 -420
rect 5850 -390 5890 -385
rect 5850 -420 5855 -390
rect 5885 -420 5890 -390
rect 5850 -425 5890 -420
rect -120 -440 -80 -435
rect -120 -470 -115 -440
rect -85 -470 -80 -440
rect -120 -475 -80 -470
rect -180 -540 -140 -535
rect -180 -570 -175 -540
rect -145 -570 -140 -540
rect -180 -575 -140 -570
rect -240 -1585 -200 -1580
rect -240 -1615 -235 -1585
rect -205 -1615 -200 -1585
rect -240 -1620 -200 -1615
rect -170 -1675 -150 -575
rect -180 -1680 -140 -1675
rect -180 -1710 -175 -1680
rect -145 -1710 -140 -1680
rect -180 -1715 -140 -1710
rect -110 -1725 -90 -475
rect -60 -490 -20 -485
rect -60 -520 -55 -490
rect -25 -520 -20 -490
rect -60 -525 -20 -520
rect -120 -1730 -80 -1725
rect -120 -1760 -115 -1730
rect -85 -1760 -80 -1730
rect -120 -1765 -80 -1760
rect -50 -1775 -30 -525
rect 1855 -870 1895 -865
rect 1855 -900 1860 -870
rect 1890 -900 1895 -870
rect 1855 -905 1895 -900
rect 1955 -925 1975 -425
rect 3805 -870 3845 -865
rect 3805 -900 3810 -870
rect 3840 -900 3845 -870
rect 3805 -905 3845 -900
rect 3910 -925 3930 -425
rect 5755 -870 5795 -865
rect 5755 -900 5760 -870
rect 5790 -900 5795 -870
rect 5755 -905 5795 -900
rect 5860 -925 5880 -425
rect 7705 -870 7745 -865
rect 7705 -900 7710 -870
rect 7740 -900 7745 -870
rect 7705 -905 7745 -900
rect 7780 -920 7820 -915
rect 7780 -925 7785 -920
rect 1895 -945 1975 -925
rect 3840 -945 3930 -925
rect 5790 -945 5880 -925
rect 7720 -945 7785 -925
rect 7780 -950 7785 -945
rect 7815 -950 7820 -920
rect 7780 -955 7820 -950
rect 1760 -1290 5880 -1270
rect 7925 -1400 7965 -1395
rect 7925 -1430 7930 -1400
rect 7960 -1430 7965 -1400
rect 7925 -1435 7965 -1430
rect 7865 -1450 7905 -1445
rect 7865 -1480 7870 -1450
rect 7900 -1480 7905 -1450
rect 7865 -1485 7905 -1480
rect 7805 -1500 7845 -1495
rect 7805 -1530 7810 -1500
rect 7840 -1530 7845 -1500
rect 7805 -1535 7845 -1530
rect 7745 -1550 7795 -1545
rect 7745 -1580 7750 -1550
rect 7780 -1580 7795 -1550
rect 7745 -1585 7795 -1580
rect 1780 -1645 5900 -1625
rect 1945 -1680 1985 -1675
rect 1945 -1710 1950 -1680
rect 1980 -1710 1985 -1680
rect 1945 -1715 1985 -1710
rect 3900 -1680 3940 -1675
rect 3900 -1710 3905 -1680
rect 3935 -1710 3940 -1680
rect 3900 -1715 3940 -1710
rect 5850 -1680 5890 -1675
rect 5850 -1710 5855 -1680
rect 5885 -1710 5890 -1680
rect 5850 -1715 5890 -1710
rect -60 -1780 -20 -1775
rect -60 -1810 -55 -1780
rect -25 -1810 -20 -1780
rect -60 -1815 -20 -1810
rect 1855 -2160 1895 -2155
rect 1855 -2190 1860 -2160
rect 1890 -2190 1895 -2160
rect 1855 -2195 1895 -2190
rect 1955 -2215 1975 -1715
rect 3800 -2160 3840 -2155
rect 3800 -2190 3805 -2160
rect 3835 -2190 3840 -2160
rect 3800 -2195 3840 -2190
rect 3910 -2215 3930 -1715
rect 5755 -2160 5795 -2155
rect 5755 -2190 5760 -2160
rect 5790 -2190 5795 -2160
rect 5755 -2195 5795 -2190
rect 5860 -2215 5880 -1715
rect 7705 -2160 7745 -2155
rect 7705 -2190 7710 -2160
rect 7740 -2190 7745 -2160
rect 7705 -2195 7745 -2190
rect 1895 -2235 1975 -2215
rect 3840 -2235 3930 -2215
rect 5795 -2235 5880 -2215
rect 7725 -2260 7745 -2215
rect 7710 -2270 7760 -2260
rect 7710 -2300 7720 -2270
rect 7750 -2300 7760 -2270
rect 7710 -2310 7760 -2300
rect 1780 -2580 5960 -2560
rect 7595 -2600 7635 -2595
rect 7595 -2605 7600 -2600
rect 420 -2625 7600 -2605
rect 420 -3000 440 -2625
rect 7595 -2630 7600 -2625
rect 7630 -2630 7635 -2600
rect 7595 -2635 7635 -2630
rect 7775 -2655 7795 -1585
rect 480 -2675 7795 -2655
rect 480 -2950 500 -2675
rect 7815 -2690 7835 -1535
rect 1590 -2710 7835 -2690
rect 1590 -2770 1610 -2710
rect 7875 -2725 7895 -1485
rect 2800 -2745 7895 -2725
rect 1580 -2775 1620 -2770
rect 1580 -2805 1585 -2775
rect 1615 -2805 1620 -2775
rect 2800 -2790 2820 -2745
rect 7935 -2760 7955 -1435
rect 7980 -2595 8000 345
rect 7970 -2600 8010 -2595
rect 7970 -2630 7975 -2600
rect 8005 -2630 8010 -2600
rect 7970 -2635 8010 -2630
rect 3985 -2780 7955 -2760
rect 1580 -2810 1620 -2805
rect 2790 -2795 2830 -2790
rect 3985 -2795 4005 -2780
rect 2790 -2825 2795 -2795
rect 2825 -2825 2830 -2795
rect 2790 -2830 2830 -2825
rect 3975 -2800 4015 -2795
rect 3975 -2830 3980 -2800
rect 4010 -2830 4015 -2800
rect 3975 -2835 4015 -2830
rect 2320 -2880 5310 -2865
rect 2320 -2885 3280 -2880
rect 3475 -2885 5310 -2880
rect 470 -2955 510 -2950
rect 470 -2985 475 -2955
rect 505 -2985 510 -2955
rect 470 -2990 510 -2985
rect 410 -3005 450 -3000
rect 410 -3035 415 -3005
rect 445 -3035 450 -3005
rect 410 -3040 450 -3035
rect 3665 -3285 3705 -3280
rect 1315 -3290 1355 -3285
rect 1315 -3320 1320 -3290
rect 1350 -3320 1355 -3290
rect 1315 -3325 1355 -3320
rect 2490 -3290 2530 -3285
rect 2490 -3320 2495 -3290
rect 2525 -3320 2530 -3290
rect 3665 -3315 3670 -3285
rect 3700 -3315 3705 -3285
rect 3665 -3320 3705 -3315
rect 4840 -3290 4880 -3285
rect 4840 -3320 4845 -3290
rect 4875 -3320 4880 -3290
rect 2490 -3325 2530 -3320
rect 4840 -3325 4880 -3320
rect 6015 -3290 6055 -3285
rect 6015 -3320 6020 -3290
rect 6050 -3320 6055 -3290
rect 6015 -3325 6055 -3320
rect 1145 -3580 5330 -3560
<< via1 >>
rect 1920 870 1950 900
rect 3870 870 3900 900
rect 5820 870 5850 900
rect 1860 390 1890 420
rect 3810 390 3840 420
rect 5760 390 5790 420
rect 7710 390 7740 420
rect -535 -75 -505 -45
rect -475 -125 -445 -95
rect -535 -1365 -505 -1335
rect -415 -175 -385 -145
rect -475 -1415 -445 -1385
rect -355 -225 -325 -195
rect -415 -1465 -385 -1435
rect -295 -275 -265 -245
rect -355 -1515 -325 -1485
rect -235 -325 -205 -295
rect -295 -1565 -265 -1535
rect 1950 -420 1980 -390
rect 3905 -420 3935 -390
rect 5855 -420 5885 -390
rect -115 -470 -85 -440
rect -175 -570 -145 -540
rect -235 -1615 -205 -1585
rect -175 -1710 -145 -1680
rect -55 -520 -25 -490
rect -115 -1760 -85 -1730
rect 1860 -900 1890 -870
rect 3810 -900 3840 -870
rect 5760 -900 5790 -870
rect 7710 -900 7740 -870
rect 7785 -950 7815 -920
rect 7930 -1430 7960 -1400
rect 7870 -1480 7900 -1450
rect 7810 -1530 7840 -1500
rect 7750 -1580 7780 -1550
rect 1950 -1710 1980 -1680
rect 3905 -1710 3935 -1680
rect 5855 -1710 5885 -1680
rect -55 -1810 -25 -1780
rect 1860 -2190 1890 -2160
rect 3805 -2190 3835 -2160
rect 5760 -2190 5790 -2160
rect 7710 -2190 7740 -2160
rect 7720 -2300 7750 -2270
rect 7600 -2630 7630 -2600
rect 1585 -2805 1615 -2775
rect 7975 -2630 8005 -2600
rect 2795 -2825 2825 -2795
rect 3980 -2830 4010 -2800
rect 475 -2985 505 -2955
rect 415 -3035 445 -3005
rect 1320 -3320 1350 -3290
rect 2495 -3320 2525 -3290
rect 3670 -3315 3700 -3285
rect 4845 -3320 4875 -3290
rect 6020 -3320 6050 -3290
<< metal2 >>
rect -620 1130 5795 1150
rect -620 1095 5755 1115
rect -620 1060 3845 1080
rect -620 1025 3805 1045
rect -620 990 1895 1010
rect -620 955 1855 975
rect -620 920 5 940
rect -620 885 -35 905
rect -620 850 -75 870
rect -95 795 -75 850
rect -55 845 -35 885
rect -15 875 5 920
rect -55 825 5 845
rect 1835 795 1855 955
rect 1875 845 1895 990
rect 1915 900 1955 905
rect 1915 870 1920 900
rect 1950 870 1955 900
rect 1915 865 1955 870
rect 1875 825 1955 845
rect 3785 795 3805 1025
rect 3825 845 3845 1060
rect 3865 900 3905 905
rect 3865 870 3870 900
rect 3900 895 3905 900
rect 3900 875 3915 895
rect 3900 870 3905 875
rect 3865 865 3905 870
rect 3825 825 3905 845
rect 5735 795 5755 1095
rect 5775 845 5795 1130
rect 5815 900 5855 905
rect 5815 870 5820 900
rect 5850 895 5855 900
rect 5850 875 5865 895
rect 5850 870 5855 875
rect 5815 865 5855 870
rect 5775 825 5860 845
rect -95 775 5 795
rect 1835 775 1955 795
rect 3785 775 3905 795
rect 5735 775 5905 795
rect 1855 420 1895 425
rect 1855 390 1860 420
rect 1890 390 1895 420
rect 1855 385 1895 390
rect 3805 420 3845 425
rect 3805 390 3810 420
rect 3840 390 3845 420
rect 3805 385 3845 390
rect 5755 420 5795 425
rect 5755 390 5760 420
rect 5790 390 5795 420
rect 5755 385 5795 390
rect 7705 420 7745 425
rect 7705 390 7710 420
rect 7740 390 7745 420
rect 7705 385 7745 390
rect -540 -45 -500 -40
rect -540 -50 -535 -45
rect -625 -70 -535 -50
rect -540 -75 -535 -70
rect -505 -50 -500 -45
rect -505 -70 1830 -50
rect -505 -75 -500 -70
rect -540 -80 -500 -75
rect -480 -95 -440 -90
rect -480 -100 -475 -95
rect -625 -120 -475 -100
rect -480 -125 -475 -120
rect -445 -100 -440 -95
rect -445 -120 1790 -100
rect -445 -125 -440 -120
rect -480 -130 -440 -125
rect -420 -145 -380 -140
rect -420 -150 -415 -145
rect -625 -170 -415 -150
rect -420 -175 -415 -170
rect -385 -150 -380 -145
rect -385 -170 1750 -150
rect -385 -175 -380 -170
rect -420 -180 -380 -175
rect -360 -195 -320 -190
rect -360 -200 -355 -195
rect -625 -220 -355 -200
rect -360 -225 -355 -220
rect -325 -200 -320 -195
rect -325 -220 1710 -200
rect -325 -225 -320 -220
rect -360 -230 -320 -225
rect -300 -245 -260 -240
rect -300 -250 -295 -245
rect -625 -270 -295 -250
rect -300 -275 -295 -270
rect -265 -250 -260 -245
rect 1690 -245 1710 -220
rect 1730 -210 1750 -170
rect 1770 -175 1790 -120
rect 1810 -140 1830 -70
rect 1865 -105 1885 385
rect 3815 -70 3835 385
rect 5765 -35 5785 385
rect 7715 0 7735 385
rect 7715 -20 7775 0
rect 5765 -55 7775 -35
rect 3815 -90 7775 -70
rect 1865 -125 7775 -105
rect 1810 -160 5795 -140
rect 1770 -195 5755 -175
rect 1730 -230 3845 -210
rect -265 -270 1670 -250
rect 1690 -265 3805 -245
rect -265 -275 -260 -270
rect -300 -280 -260 -275
rect 1650 -280 1670 -270
rect -240 -295 -200 -290
rect -240 -300 -235 -295
rect -625 -320 -235 -300
rect -240 -325 -235 -320
rect -205 -300 -200 -295
rect 1650 -300 1895 -280
rect -205 -315 1630 -300
rect -205 -320 1855 -315
rect -205 -325 -200 -320
rect -240 -330 -200 -325
rect 1610 -335 1855 -320
rect -625 -415 5 -395
rect -120 -440 -80 -435
rect -120 -445 -115 -440
rect -625 -465 -115 -445
rect -120 -470 -115 -465
rect -85 -445 -80 -440
rect -85 -465 5 -445
rect -85 -470 -80 -465
rect -120 -475 -80 -470
rect -60 -490 -20 -485
rect -60 -495 -55 -490
rect -625 -515 -55 -495
rect -60 -520 -55 -515
rect -25 -495 -20 -490
rect 1835 -495 1855 -335
rect 1875 -445 1895 -300
rect 1945 -390 1985 -385
rect 1945 -420 1950 -390
rect 1980 -420 1985 -390
rect 1945 -425 1985 -420
rect 1875 -465 1955 -445
rect 3785 -495 3805 -265
rect 3825 -445 3845 -230
rect 3900 -390 3940 -385
rect 3900 -420 3905 -390
rect 3935 -420 3940 -390
rect 3900 -425 3940 -420
rect 3825 -465 3920 -445
rect 5735 -495 5755 -195
rect 5775 -445 5795 -160
rect 5850 -390 5890 -385
rect 5850 -420 5855 -390
rect 5885 -420 5890 -390
rect 5850 -425 5890 -420
rect 5775 -465 5870 -445
rect -25 -515 5 -495
rect 1835 -515 1950 -495
rect 3785 -515 3905 -495
rect 5735 -515 5885 -495
rect -25 -520 -20 -515
rect -60 -525 -20 -520
rect -180 -540 -140 -535
rect -180 -545 -175 -540
rect -625 -565 -175 -545
rect -180 -570 -175 -565
rect -145 -570 -140 -540
rect -180 -575 -140 -570
rect 1855 -870 1895 -865
rect 1855 -900 1860 -870
rect 1890 -900 1895 -870
rect 1855 -905 1895 -900
rect 3805 -870 3845 -865
rect 3805 -900 3810 -870
rect 3840 -900 3845 -870
rect 3805 -905 3845 -900
rect 5755 -870 5795 -865
rect 5755 -900 5760 -870
rect 5790 -900 5795 -870
rect 5755 -905 5795 -900
rect 7705 -870 7745 -865
rect 7705 -900 7710 -870
rect 7740 -900 7745 -870
rect 7705 -905 7745 -900
rect -540 -1335 -500 -1330
rect -540 -1365 -535 -1335
rect -505 -1340 -500 -1335
rect -505 -1360 1830 -1340
rect -505 -1365 -500 -1360
rect -540 -1370 -500 -1365
rect -480 -1385 -440 -1380
rect -480 -1415 -475 -1385
rect -445 -1390 -440 -1385
rect -445 -1410 1790 -1390
rect -445 -1415 -440 -1410
rect -480 -1420 -440 -1415
rect -420 -1435 -380 -1430
rect -420 -1465 -415 -1435
rect -385 -1440 -380 -1435
rect -385 -1460 1750 -1440
rect -385 -1465 -380 -1460
rect -420 -1470 -380 -1465
rect -360 -1485 -320 -1480
rect -360 -1515 -355 -1485
rect -325 -1490 -320 -1485
rect -325 -1510 1710 -1490
rect -325 -1515 -320 -1510
rect -360 -1520 -320 -1515
rect -300 -1535 -260 -1530
rect -300 -1565 -295 -1535
rect -265 -1540 -260 -1535
rect 1690 -1535 1710 -1510
rect 1730 -1500 1750 -1460
rect 1770 -1465 1790 -1410
rect 1810 -1430 1830 -1360
rect 1865 -1395 1885 -905
rect 3815 -1360 3835 -905
rect 5765 -1325 5785 -905
rect 5765 -1345 7490 -1325
rect 3815 -1380 7440 -1360
rect 1865 -1415 7390 -1395
rect 1810 -1450 5795 -1430
rect 1770 -1485 5755 -1465
rect 1730 -1520 3845 -1500
rect -265 -1560 1670 -1540
rect 1690 -1555 3805 -1535
rect -265 -1565 -260 -1560
rect -300 -1570 -260 -1565
rect 1650 -1570 1670 -1560
rect -240 -1585 -200 -1580
rect -240 -1615 -235 -1585
rect -205 -1590 -200 -1585
rect 1650 -1590 1895 -1570
rect -205 -1605 1630 -1590
rect -205 -1610 1855 -1605
rect -205 -1615 -200 -1610
rect -240 -1620 -200 -1615
rect 1610 -1625 1855 -1610
rect -180 -1680 -140 -1675
rect -180 -1710 -175 -1680
rect -145 -1685 -140 -1680
rect -145 -1705 5 -1685
rect -145 -1710 -140 -1705
rect -180 -1715 -140 -1710
rect -120 -1730 -80 -1725
rect -120 -1760 -115 -1730
rect -85 -1735 -80 -1730
rect -85 -1755 5 -1735
rect -85 -1760 -80 -1755
rect -120 -1765 -80 -1760
rect -60 -1780 -20 -1775
rect -60 -1810 -55 -1780
rect -25 -1785 -20 -1780
rect 1835 -1785 1855 -1625
rect 1875 -1735 1895 -1590
rect 1945 -1680 1985 -1675
rect 1945 -1710 1950 -1680
rect 1980 -1710 1985 -1680
rect 1945 -1715 1985 -1710
rect 1875 -1755 1950 -1735
rect 3785 -1785 3805 -1555
rect 3825 -1735 3845 -1520
rect 3900 -1680 3940 -1675
rect 3900 -1710 3905 -1680
rect 3935 -1710 3940 -1680
rect 3900 -1715 3940 -1710
rect 3825 -1755 3905 -1735
rect 5735 -1785 5755 -1485
rect 5775 -1735 5795 -1450
rect 7370 -1555 7390 -1415
rect 7420 -1505 7440 -1380
rect 7470 -1455 7490 -1345
rect 7715 -1405 7735 -905
rect 7780 -920 7820 -915
rect 7780 -950 7785 -920
rect 7815 -925 7820 -920
rect 7815 -945 8095 -925
rect 7815 -950 7820 -945
rect 7780 -955 7820 -950
rect 7925 -1400 7965 -1395
rect 7925 -1405 7930 -1400
rect 7715 -1425 7930 -1405
rect 7925 -1430 7930 -1425
rect 7960 -1430 7965 -1400
rect 7925 -1435 7965 -1430
rect 7865 -1450 7905 -1445
rect 7865 -1455 7870 -1450
rect 7470 -1475 7870 -1455
rect 7865 -1480 7870 -1475
rect 7900 -1480 7905 -1450
rect 7865 -1485 7905 -1480
rect 7805 -1500 7845 -1495
rect 7805 -1505 7810 -1500
rect 7420 -1525 7810 -1505
rect 7805 -1530 7810 -1525
rect 7840 -1530 7845 -1500
rect 7805 -1535 7845 -1530
rect 7745 -1550 7795 -1545
rect 7745 -1555 7750 -1550
rect 7370 -1575 7750 -1555
rect 7745 -1580 7750 -1575
rect 7780 -1580 7795 -1550
rect 7745 -1585 7795 -1580
rect 5850 -1680 5890 -1675
rect 5850 -1710 5855 -1680
rect 5885 -1710 5890 -1680
rect 5850 -1715 5890 -1710
rect 5775 -1755 5910 -1735
rect -25 -1805 5 -1785
rect 1835 -1805 1950 -1785
rect 3785 -1805 3905 -1785
rect 5735 -1805 5855 -1785
rect -25 -1810 -20 -1805
rect -60 -1815 -20 -1810
rect 1855 -2160 1895 -2155
rect 1855 -2190 1860 -2160
rect 1890 -2190 1895 -2160
rect 1855 -2195 1895 -2190
rect 3800 -2160 3840 -2155
rect 3800 -2190 3805 -2160
rect 3835 -2190 3840 -2160
rect 3800 -2195 3840 -2190
rect 5755 -2160 5795 -2155
rect 5755 -2190 5760 -2160
rect 5790 -2190 5795 -2160
rect 5755 -2195 5795 -2190
rect 7705 -2160 7745 -2155
rect 7705 -2190 7710 -2160
rect 7740 -2165 7745 -2160
rect 7740 -2185 8060 -2165
rect 7740 -2190 7745 -2185
rect 7705 -2195 7745 -2190
rect 1865 -2675 1885 -2195
rect 520 -2695 1885 -2675
rect 520 -2910 540 -2695
rect 3810 -2710 3830 -2195
rect 1700 -2730 3830 -2710
rect 1580 -2775 1620 -2770
rect 1580 -2805 1585 -2775
rect 1615 -2805 1620 -2775
rect 1580 -2810 1620 -2805
rect 520 -2930 610 -2910
rect 470 -2955 510 -2950
rect 470 -2985 475 -2955
rect 505 -2960 510 -2955
rect 1590 -2960 1610 -2810
rect 1700 -2910 1720 -2730
rect 5765 -2750 5785 -2195
rect 7710 -2270 7760 -2260
rect 7710 -2300 7720 -2270
rect 7750 -2300 7760 -2270
rect 7710 -2310 7760 -2300
rect 7595 -2600 7635 -2595
rect 7595 -2630 7600 -2600
rect 7630 -2605 7635 -2600
rect 7970 -2600 8010 -2595
rect 7970 -2605 7975 -2600
rect 7630 -2625 7975 -2605
rect 7630 -2630 7635 -2625
rect 7595 -2635 7635 -2630
rect 7970 -2630 7975 -2625
rect 8005 -2630 8010 -2600
rect 7970 -2635 8010 -2630
rect 2850 -2770 5785 -2750
rect 2790 -2795 2830 -2790
rect 2790 -2825 2795 -2795
rect 2825 -2825 2830 -2795
rect 2790 -2830 2830 -2825
rect 1700 -2930 1785 -2910
rect 2800 -2955 2820 -2830
rect 2850 -2905 2870 -2770
rect 8040 -2790 8060 -2185
rect 3975 -2800 4015 -2795
rect 3975 -2830 3980 -2800
rect 4010 -2830 4015 -2800
rect 3975 -2835 4015 -2830
rect 4055 -2810 8060 -2790
rect 2850 -2925 2960 -2905
rect 505 -2980 615 -2960
rect 505 -2985 510 -2980
rect 470 -2990 510 -2985
rect 1010 -2990 1485 -2970
rect 1590 -2980 1785 -2960
rect 410 -3005 450 -3000
rect 410 -3035 415 -3005
rect 445 -3010 450 -3005
rect 1010 -3010 1030 -2990
rect 445 -3030 610 -3010
rect 980 -3030 1030 -3010
rect 1465 -3010 1485 -2990
rect 2190 -2985 2610 -2965
rect 2800 -2975 2960 -2955
rect 3985 -2960 4005 -2835
rect 4055 -2910 4075 -2810
rect 8075 -2825 8095 -945
rect 5115 -2845 8095 -2825
rect 4055 -2930 4135 -2910
rect 5115 -2960 5135 -2845
rect 5260 -2870 5930 -2860
rect 7710 -2870 7760 -2865
rect 5260 -2880 7715 -2870
rect 5260 -2910 5280 -2880
rect 5910 -2890 7715 -2880
rect 7710 -2910 7715 -2890
rect 7755 -2910 7760 -2870
rect 5260 -2930 5390 -2910
rect 7710 -2915 7760 -2910
rect 2190 -3010 2210 -2985
rect 1465 -3030 1795 -3010
rect 2165 -3030 2210 -3010
rect 2590 -3005 2610 -2985
rect 3365 -2980 3790 -2960
rect 3985 -2980 4135 -2960
rect 4540 -2980 4905 -2960
rect 5115 -2980 5310 -2960
rect 3365 -3005 3385 -2980
rect 2590 -3025 2960 -3005
rect 3340 -3025 3385 -3005
rect 3770 -3010 3790 -2980
rect 4540 -3010 4560 -2980
rect 3770 -3030 4135 -3010
rect 4490 -3030 4560 -3010
rect 4885 -3010 4905 -2980
rect 4885 -3030 5310 -3010
rect 445 -3035 450 -3030
rect 410 -3040 450 -3035
rect 3665 -3285 3705 -3280
rect 1315 -3290 1355 -3285
rect 1315 -3320 1320 -3290
rect 1350 -3320 1355 -3290
rect 1315 -3325 1355 -3320
rect 2490 -3290 2530 -3285
rect 2490 -3320 2495 -3290
rect 2525 -3320 2530 -3290
rect 3665 -3315 3670 -3285
rect 3700 -3315 3705 -3285
rect 3665 -3320 3705 -3315
rect 4840 -3290 4880 -3285
rect 4840 -3320 4845 -3290
rect 4875 -3320 4880 -3290
rect 2490 -3325 2530 -3320
rect 1325 -3630 1345 -3325
rect 2500 -3595 2520 -3325
rect 3675 -3560 3695 -3320
rect 4840 -3325 4880 -3320
rect 6015 -3290 6055 -3285
rect 6015 -3320 6020 -3290
rect 6050 -3295 6055 -3290
rect 6050 -3315 7790 -3295
rect 6050 -3320 6055 -3315
rect 6015 -3325 6055 -3320
rect 4850 -3525 4870 -3325
rect 6200 -3350 7790 -3330
rect 6200 -3525 6220 -3350
rect 4850 -3545 6220 -3525
rect 6240 -3385 7790 -3365
rect 6240 -3560 6260 -3385
rect 3675 -3580 6260 -3560
rect 6280 -3420 7790 -3400
rect 6280 -3595 6300 -3420
rect 2500 -3615 6300 -3595
rect 6320 -3455 7790 -3435
rect 6320 -3630 6340 -3455
rect 1325 -3650 6340 -3630
<< via2 >>
rect 7720 -2300 7750 -2270
rect 7715 -2910 7755 -2870
<< metal3 >>
rect 7710 -2270 7760 -2260
rect 7710 -2300 7720 -2270
rect 7750 -2300 7760 -2270
rect 7710 -2310 7760 -2300
rect 7720 -2865 7750 -2310
rect 7710 -2870 7760 -2865
rect 7710 -2910 7715 -2870
rect 7755 -2910 7760 -2870
rect 7710 -2915 7760 -2910
use full_adder  full_adder_0
timestamp 1720452554
transform 1 0 2040 0 1 460
box -90 -460 1805 495
use full_adder  full_adder_1
timestamp 1720452554
transform 1 0 90 0 1 460
box -90 -460 1805 495
use full_adder  full_adder_2
timestamp 1720452554
transform 1 0 3990 0 1 460
box -90 -460 1805 495
use full_adder  full_adder_3
timestamp 1720452554
transform 1 0 5940 0 1 -830
box -90 -460 1805 495
use full_adder  full_adder_4
timestamp 1720452554
transform 1 0 5940 0 1 460
box -90 -460 1805 495
use full_adder  full_adder_5
timestamp 1720452554
transform 1 0 90 0 1 -830
box -90 -460 1805 495
use full_adder  full_adder_6
timestamp 1720452554
transform 1 0 2035 0 1 -830
box -90 -460 1805 495
use full_adder  full_adder_7
timestamp 1720452554
transform 1 0 3990 0 1 -830
box -90 -460 1805 495
use full_adder  full_adder_8
timestamp 1720452554
transform 1 0 2035 0 1 -2120
box -90 -460 1805 495
use full_adder  full_adder_9
timestamp 1720452554
transform 1 0 90 0 1 -2120
box -90 -460 1805 495
use full_adder  full_adder_10
timestamp 1720452554
transform 1 0 3990 0 1 -2120
box -90 -460 1805 495
use full_adder  full_adder_11
timestamp 1720452554
transform 1 0 5940 0 1 -2120
box -90 -460 1805 495
use mux_2to1  mux_2to1_0
timestamp 1720464950
transform 1 0 -505 0 1 -3705
box 1115 125 1820 840
use mux_2to1  mux_2to1_1
timestamp 1720464950
transform 1 0 670 0 1 -3705
box 1115 125 1820 840
use mux_2to1  mux_2to1_2
timestamp 1720464950
transform 1 0 1845 0 1 -3700
box 1115 125 1820 840
use mux_2to1  mux_2to1_3
timestamp 1720464950
transform 1 0 3020 0 1 -3705
box 1115 125 1820 840
use mux_2to1  mux_2to1_4
timestamp 1720464950
transform 1 0 4195 0 1 -3705
box 1115 125 1820 840
<< labels >>
rlabel metal2 7760 -125 7770 -105 1 s0
rlabel metal2 7760 -90 7770 -70 1 s1
rlabel metal2 7760 -55 7770 -35 1 s2
rlabel metal2 7760 -20 7770 0 1 s3
rlabel metal2 7775 -3315 7785 -3295 1 cout
rlabel metal2 7775 -3455 7785 -3435 1 s4
rlabel metal2 7775 -3420 7785 -3400 1 s5
rlabel metal2 7775 -3385 7785 -3365 1 s6
rlabel metal2 7775 -3350 7785 -3330 1 s7
rlabel metal2 -610 850 -600 870 1 a0
rlabel metal2 -610 885 -600 905 1 b0
rlabel metal2 -610 955 -600 975 1 a1
rlabel metal2 -610 1025 -600 1045 1 a2
rlabel metal2 -610 1095 -600 1115 1 a3
rlabel metal2 -610 990 -600 1010 1 b1
rlabel metal2 -610 1060 -600 1080 1 b2
rlabel metal2 -610 1130 -600 1150 1 b3
rlabel metal2 -615 -415 -605 -395 1 cin0
rlabel metal2 -615 -515 -605 -495 1 a4
rlabel metal2 -615 -320 -605 -300 1 a5
rlabel metal2 -615 -220 -605 -200 1 a6
rlabel metal2 -615 -120 -605 -100 1 a7
rlabel metal2 -615 -465 -605 -445 1 b4
rlabel metal2 -615 -270 -605 -250 1 b5
rlabel metal2 -615 -170 -605 -150 1 b6
rlabel metal2 -615 -70 -605 -50 1 b7
rlabel metal2 -615 -565 -605 -545 1 cin1
rlabel metal1 1395 -3570 1395 -3570 1 gnd
rlabel metal1 2610 -2875 2610 -2875 1 vdd
rlabel metal1 1820 -2575 1820 -2575 1 gnd
rlabel metal1 1805 -1635 1805 -1635 1 vdd
rlabel metal1 1815 -1285 1815 -1285 1 gnd
rlabel metal1 1805 -350 1805 -350 1 vdd
rlabel metal1 1820 5 1820 5 1 gnd
rlabel metal1 1915 940 1915 940 1 vdd
rlabel metal2 -610 920 -600 940 1 cin0
<< end >>
